`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Mul(
  input  [1:0] io_in0,
  input  [1:0] io_in1,
  output [1:0] io_out
);
  wire [3:0] _T_5;
  assign _T_5 = io_in0 * io_in1;
  assign io_out = _T_5[1:0];
endmodule
module VectorElemAdd(
  input  [1:0] io_input_0,
  input  [1:0] io_input_1,
  input  [1:0] io_input_2,
  input  [1:0] io_input_3,
  input  [1:0] io_input_4,
  input  [1:0] io_input_5,
  input  [1:0] io_input_6,
  input  [1:0] io_input_7,
  input  [1:0] io_input_8,
  output [1:0] io_out
);
  wire [2:0] _T_17;
  wire [1:0] _T_18;
  wire [2:0] _T_19;
  wire [1:0] _T_20;
  wire [2:0] _T_21;
  wire [1:0] _T_22;
  wire [2:0] _T_23;
  wire [1:0] _T_24;
  wire [2:0] _T_25;
  wire [1:0] _T_26;
  wire [2:0] _T_27;
  wire [1:0] _T_28;
  wire [2:0] _T_29;
  wire [1:0] _T_30;
  wire [2:0] _T_31;
  wire [1:0] _T_32;
  assign _T_17 = io_input_0 + io_input_1;
  assign _T_18 = _T_17[1:0];
  assign _T_19 = _T_18 + io_input_2;
  assign _T_20 = _T_19[1:0];
  assign _T_21 = _T_20 + io_input_3;
  assign _T_22 = _T_21[1:0];
  assign _T_23 = _T_22 + io_input_4;
  assign _T_24 = _T_23[1:0];
  assign _T_25 = _T_24 + io_input_5;
  assign _T_26 = _T_25[1:0];
  assign _T_27 = _T_26 + io_input_6;
  assign _T_28 = _T_27[1:0];
  assign _T_29 = _T_28 + io_input_7;
  assign _T_30 = _T_29[1:0];
  assign _T_31 = _T_30 + io_input_8;
  assign _T_32 = _T_31[1:0];
  assign io_out = _T_32;
endmodule
module VectorMul(
  input        clock,
  input        reset,
  input  [1:0] io_vec1_0,
  input  [1:0] io_vec1_1,
  input  [1:0] io_vec1_2,
  input  [1:0] io_vec1_3,
  input  [1:0] io_vec1_4,
  input  [1:0] io_vec1_5,
  input  [1:0] io_vec1_6,
  input  [1:0] io_vec1_7,
  input  [1:0] io_vec1_8,
  input  [1:0] io_vec2_0,
  input  [1:0] io_vec2_1,
  input  [1:0] io_vec2_2,
  input  [1:0] io_vec2_3,
  input  [1:0] io_vec2_4,
  input  [1:0] io_vec2_5,
  input  [1:0] io_vec2_6,
  input  [1:0] io_vec2_7,
  input  [1:0] io_vec2_8,
  output [1:0] io_out
);
  wire [1:0] Mul_io_in0;
  wire [1:0] Mul_io_in1;
  wire [1:0] Mul_io_out;
  wire [1:0] Mul_1_io_in0;
  wire [1:0] Mul_1_io_in1;
  wire [1:0] Mul_1_io_out;
  wire [1:0] Mul_2_io_in0;
  wire [1:0] Mul_2_io_in1;
  wire [1:0] Mul_2_io_out;
  wire [1:0] Mul_3_io_in0;
  wire [1:0] Mul_3_io_in1;
  wire [1:0] Mul_3_io_out;
  wire [1:0] Mul_4_io_in0;
  wire [1:0] Mul_4_io_in1;
  wire [1:0] Mul_4_io_out;
  wire [1:0] Mul_5_io_in0;
  wire [1:0] Mul_5_io_in1;
  wire [1:0] Mul_5_io_out;
  wire [1:0] Mul_6_io_in0;
  wire [1:0] Mul_6_io_in1;
  wire [1:0] Mul_6_io_out;
  wire [1:0] Mul_7_io_in0;
  wire [1:0] Mul_7_io_in1;
  wire [1:0] Mul_7_io_out;
  wire [1:0] Mul_8_io_in0;
  wire [1:0] Mul_8_io_in1;
  wire [1:0] Mul_8_io_out;
  reg [1:0] quotient_0;
  reg [31:0] _RAND_0;
  reg [1:0] quotient_1;
  reg [31:0] _RAND_1;
  reg [1:0] quotient_2;
  reg [31:0] _RAND_2;
  reg [1:0] quotient_3;
  reg [31:0] _RAND_3;
  reg [1:0] quotient_4;
  reg [31:0] _RAND_4;
  reg [1:0] quotient_5;
  reg [31:0] _RAND_5;
  reg [1:0] quotient_6;
  reg [31:0] _RAND_6;
  reg [1:0] quotient_7;
  reg [31:0] _RAND_7;
  reg [1:0] quotient_8;
  reg [31:0] _RAND_8;
  wire [1:0] VectorElemAdd_io_input_0;
  wire [1:0] VectorElemAdd_io_input_1;
  wire [1:0] VectorElemAdd_io_input_2;
  wire [1:0] VectorElemAdd_io_input_3;
  wire [1:0] VectorElemAdd_io_input_4;
  wire [1:0] VectorElemAdd_io_input_5;
  wire [1:0] VectorElemAdd_io_input_6;
  wire [1:0] VectorElemAdd_io_input_7;
  wire [1:0] VectorElemAdd_io_input_8;
  wire [1:0] VectorElemAdd_io_out;
  Mul Mul (
    .io_in0(Mul_io_in0),
    .io_in1(Mul_io_in1),
    .io_out(Mul_io_out)
  );
  Mul Mul_1 (
    .io_in0(Mul_1_io_in0),
    .io_in1(Mul_1_io_in1),
    .io_out(Mul_1_io_out)
  );
  Mul Mul_2 (
    .io_in0(Mul_2_io_in0),
    .io_in1(Mul_2_io_in1),
    .io_out(Mul_2_io_out)
  );
  Mul Mul_3 (
    .io_in0(Mul_3_io_in0),
    .io_in1(Mul_3_io_in1),
    .io_out(Mul_3_io_out)
  );
  Mul Mul_4 (
    .io_in0(Mul_4_io_in0),
    .io_in1(Mul_4_io_in1),
    .io_out(Mul_4_io_out)
  );
  Mul Mul_5 (
    .io_in0(Mul_5_io_in0),
    .io_in1(Mul_5_io_in1),
    .io_out(Mul_5_io_out)
  );
  Mul Mul_6 (
    .io_in0(Mul_6_io_in0),
    .io_in1(Mul_6_io_in1),
    .io_out(Mul_6_io_out)
  );
  Mul Mul_7 (
    .io_in0(Mul_7_io_in0),
    .io_in1(Mul_7_io_in1),
    .io_out(Mul_7_io_out)
  );
  Mul Mul_8 (
    .io_in0(Mul_8_io_in0),
    .io_in1(Mul_8_io_in1),
    .io_out(Mul_8_io_out)
  );
  VectorElemAdd VectorElemAdd (
    .io_input_0(VectorElemAdd_io_input_0),
    .io_input_1(VectorElemAdd_io_input_1),
    .io_input_2(VectorElemAdd_io_input_2),
    .io_input_3(VectorElemAdd_io_input_3),
    .io_input_4(VectorElemAdd_io_input_4),
    .io_input_5(VectorElemAdd_io_input_5),
    .io_input_6(VectorElemAdd_io_input_6),
    .io_input_7(VectorElemAdd_io_input_7),
    .io_input_8(VectorElemAdd_io_input_8),
    .io_out(VectorElemAdd_io_out)
  );
  assign io_out = VectorElemAdd_io_out;
  assign Mul_io_in0 = io_vec1_0;
  assign Mul_io_in1 = io_vec2_0;
  assign Mul_1_io_in0 = io_vec1_1;
  assign Mul_1_io_in1 = io_vec2_1;
  assign Mul_2_io_in0 = io_vec1_2;
  assign Mul_2_io_in1 = io_vec2_2;
  assign Mul_3_io_in0 = io_vec1_3;
  assign Mul_3_io_in1 = io_vec2_3;
  assign Mul_4_io_in0 = io_vec1_4;
  assign Mul_4_io_in1 = io_vec2_4;
  assign Mul_5_io_in0 = io_vec1_5;
  assign Mul_5_io_in1 = io_vec2_5;
  assign Mul_6_io_in0 = io_vec1_6;
  assign Mul_6_io_in1 = io_vec2_6;
  assign Mul_7_io_in0 = io_vec1_7;
  assign Mul_7_io_in1 = io_vec2_7;
  assign Mul_8_io_in0 = io_vec1_8;
  assign Mul_8_io_in1 = io_vec2_8;
  assign VectorElemAdd_io_input_0 = quotient_0;
  assign VectorElemAdd_io_input_1 = quotient_1;
  assign VectorElemAdd_io_input_2 = quotient_2;
  assign VectorElemAdd_io_input_3 = quotient_3;
  assign VectorElemAdd_io_input_4 = quotient_4;
  assign VectorElemAdd_io_input_5 = quotient_5;
  assign VectorElemAdd_io_input_6 = quotient_6;
  assign VectorElemAdd_io_input_7 = quotient_7;
  assign VectorElemAdd_io_input_8 = quotient_8;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  quotient_0 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  quotient_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  quotient_2 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  quotient_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  quotient_4 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  quotient_5 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  quotient_6 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  quotient_7 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  quotient_8 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      quotient_0 <= 2'h0;
    end else begin
      quotient_0 <= Mul_io_out;
    end
    if (reset) begin
      quotient_1 <= 2'h0;
    end else begin
      quotient_1 <= Mul_1_io_out;
    end
    if (reset) begin
      quotient_2 <= 2'h0;
    end else begin
      quotient_2 <= Mul_2_io_out;
    end
    if (reset) begin
      quotient_3 <= 2'h0;
    end else begin
      quotient_3 <= Mul_3_io_out;
    end
    if (reset) begin
      quotient_4 <= 2'h0;
    end else begin
      quotient_4 <= Mul_4_io_out;
    end
    if (reset) begin
      quotient_5 <= 2'h0;
    end else begin
      quotient_5 <= Mul_5_io_out;
    end
    if (reset) begin
      quotient_6 <= 2'h0;
    end else begin
      quotient_6 <= Mul_6_io_out;
    end
    if (reset) begin
      quotient_7 <= 2'h0;
    end else begin
      quotient_7 <= Mul_7_io_out;
    end
    if (reset) begin
      quotient_8 <= 2'h0;
    end else begin
      quotient_8 <= Mul_8_io_out;
    end
  end
endmodule
module Conv(
  input        clock,
  input        reset,
  input  [1:0] io_mask_0,
  input  [1:0] io_mask_1,
  input  [1:0] io_mask_2,
  input  [1:0] io_mask_3,
  input  [1:0] io_mask_4,
  input  [1:0] io_mask_5,
  input  [1:0] io_mask_6,
  input  [1:0] io_mask_7,
  input  [1:0] io_mask_8,
  input  [1:0] io_mask_9,
  input  [1:0] io_mask_10,
  input  [1:0] io_mask_11,
  input  [1:0] io_mask_12,
  input  [1:0] io_mask_13,
  input  [1:0] io_mask_14,
  input  [1:0] io_mask_15,
  input  [1:0] io_mask_16,
  input  [1:0] io_mask_17,
  input  [1:0] io_mask_18,
  input  [1:0] io_mask_19,
  input  [1:0] io_mask_20,
  input  [1:0] io_mask_21,
  input  [1:0] io_mask_22,
  input  [1:0] io_mask_23,
  input  [1:0] io_mask_24,
  input  [1:0] io_weights_0,
  input  [1:0] io_weights_1,
  input  [1:0] io_weights_2,
  input  [1:0] io_weights_3,
  input  [1:0] io_weights_4,
  input  [1:0] io_weights_5,
  input  [1:0] io_weights_6,
  input  [1:0] io_weights_7,
  input  [1:0] io_weights_8,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14,
  output [3:0] io_out_15,
  output [3:0] io_out_16,
  output [3:0] io_out_17,
  output [3:0] io_out_18,
  output [3:0] io_out_19,
  output [3:0] io_out_20,
  output [3:0] io_out_21,
  output [3:0] io_out_22,
  output [3:0] io_out_23,
  output [3:0] io_out_24
);
  wire  VectorMul_clock;
  wire  VectorMul_reset;
  wire [1:0] VectorMul_io_vec1_0;
  wire [1:0] VectorMul_io_vec1_1;
  wire [1:0] VectorMul_io_vec1_2;
  wire [1:0] VectorMul_io_vec1_3;
  wire [1:0] VectorMul_io_vec1_4;
  wire [1:0] VectorMul_io_vec1_5;
  wire [1:0] VectorMul_io_vec1_6;
  wire [1:0] VectorMul_io_vec1_7;
  wire [1:0] VectorMul_io_vec1_8;
  wire [1:0] VectorMul_io_vec2_0;
  wire [1:0] VectorMul_io_vec2_1;
  wire [1:0] VectorMul_io_vec2_2;
  wire [1:0] VectorMul_io_vec2_3;
  wire [1:0] VectorMul_io_vec2_4;
  wire [1:0] VectorMul_io_vec2_5;
  wire [1:0] VectorMul_io_vec2_6;
  wire [1:0] VectorMul_io_vec2_7;
  wire [1:0] VectorMul_io_vec2_8;
  wire [1:0] VectorMul_io_out;
  wire  VectorMul_1_clock;
  wire  VectorMul_1_reset;
  wire [1:0] VectorMul_1_io_vec1_0;
  wire [1:0] VectorMul_1_io_vec1_1;
  wire [1:0] VectorMul_1_io_vec1_2;
  wire [1:0] VectorMul_1_io_vec1_3;
  wire [1:0] VectorMul_1_io_vec1_4;
  wire [1:0] VectorMul_1_io_vec1_5;
  wire [1:0] VectorMul_1_io_vec1_6;
  wire [1:0] VectorMul_1_io_vec1_7;
  wire [1:0] VectorMul_1_io_vec1_8;
  wire [1:0] VectorMul_1_io_vec2_0;
  wire [1:0] VectorMul_1_io_vec2_1;
  wire [1:0] VectorMul_1_io_vec2_2;
  wire [1:0] VectorMul_1_io_vec2_3;
  wire [1:0] VectorMul_1_io_vec2_4;
  wire [1:0] VectorMul_1_io_vec2_5;
  wire [1:0] VectorMul_1_io_vec2_6;
  wire [1:0] VectorMul_1_io_vec2_7;
  wire [1:0] VectorMul_1_io_vec2_8;
  wire [1:0] VectorMul_1_io_out;
  wire  VectorMul_2_clock;
  wire  VectorMul_2_reset;
  wire [1:0] VectorMul_2_io_vec1_0;
  wire [1:0] VectorMul_2_io_vec1_1;
  wire [1:0] VectorMul_2_io_vec1_2;
  wire [1:0] VectorMul_2_io_vec1_3;
  wire [1:0] VectorMul_2_io_vec1_4;
  wire [1:0] VectorMul_2_io_vec1_5;
  wire [1:0] VectorMul_2_io_vec1_6;
  wire [1:0] VectorMul_2_io_vec1_7;
  wire [1:0] VectorMul_2_io_vec1_8;
  wire [1:0] VectorMul_2_io_vec2_0;
  wire [1:0] VectorMul_2_io_vec2_1;
  wire [1:0] VectorMul_2_io_vec2_2;
  wire [1:0] VectorMul_2_io_vec2_3;
  wire [1:0] VectorMul_2_io_vec2_4;
  wire [1:0] VectorMul_2_io_vec2_5;
  wire [1:0] VectorMul_2_io_vec2_6;
  wire [1:0] VectorMul_2_io_vec2_7;
  wire [1:0] VectorMul_2_io_vec2_8;
  wire [1:0] VectorMul_2_io_out;
  wire  VectorMul_3_clock;
  wire  VectorMul_3_reset;
  wire [1:0] VectorMul_3_io_vec1_0;
  wire [1:0] VectorMul_3_io_vec1_1;
  wire [1:0] VectorMul_3_io_vec1_2;
  wire [1:0] VectorMul_3_io_vec1_3;
  wire [1:0] VectorMul_3_io_vec1_4;
  wire [1:0] VectorMul_3_io_vec1_5;
  wire [1:0] VectorMul_3_io_vec1_6;
  wire [1:0] VectorMul_3_io_vec1_7;
  wire [1:0] VectorMul_3_io_vec1_8;
  wire [1:0] VectorMul_3_io_vec2_0;
  wire [1:0] VectorMul_3_io_vec2_1;
  wire [1:0] VectorMul_3_io_vec2_2;
  wire [1:0] VectorMul_3_io_vec2_3;
  wire [1:0] VectorMul_3_io_vec2_4;
  wire [1:0] VectorMul_3_io_vec2_5;
  wire [1:0] VectorMul_3_io_vec2_6;
  wire [1:0] VectorMul_3_io_vec2_7;
  wire [1:0] VectorMul_3_io_vec2_8;
  wire [1:0] VectorMul_3_io_out;
  wire  VectorMul_4_clock;
  wire  VectorMul_4_reset;
  wire [1:0] VectorMul_4_io_vec1_0;
  wire [1:0] VectorMul_4_io_vec1_1;
  wire [1:0] VectorMul_4_io_vec1_2;
  wire [1:0] VectorMul_4_io_vec1_3;
  wire [1:0] VectorMul_4_io_vec1_4;
  wire [1:0] VectorMul_4_io_vec1_5;
  wire [1:0] VectorMul_4_io_vec1_6;
  wire [1:0] VectorMul_4_io_vec1_7;
  wire [1:0] VectorMul_4_io_vec1_8;
  wire [1:0] VectorMul_4_io_vec2_0;
  wire [1:0] VectorMul_4_io_vec2_1;
  wire [1:0] VectorMul_4_io_vec2_2;
  wire [1:0] VectorMul_4_io_vec2_3;
  wire [1:0] VectorMul_4_io_vec2_4;
  wire [1:0] VectorMul_4_io_vec2_5;
  wire [1:0] VectorMul_4_io_vec2_6;
  wire [1:0] VectorMul_4_io_vec2_7;
  wire [1:0] VectorMul_4_io_vec2_8;
  wire [1:0] VectorMul_4_io_out;
  wire  VectorMul_5_clock;
  wire  VectorMul_5_reset;
  wire [1:0] VectorMul_5_io_vec1_0;
  wire [1:0] VectorMul_5_io_vec1_1;
  wire [1:0] VectorMul_5_io_vec1_2;
  wire [1:0] VectorMul_5_io_vec1_3;
  wire [1:0] VectorMul_5_io_vec1_4;
  wire [1:0] VectorMul_5_io_vec1_5;
  wire [1:0] VectorMul_5_io_vec1_6;
  wire [1:0] VectorMul_5_io_vec1_7;
  wire [1:0] VectorMul_5_io_vec1_8;
  wire [1:0] VectorMul_5_io_vec2_0;
  wire [1:0] VectorMul_5_io_vec2_1;
  wire [1:0] VectorMul_5_io_vec2_2;
  wire [1:0] VectorMul_5_io_vec2_3;
  wire [1:0] VectorMul_5_io_vec2_4;
  wire [1:0] VectorMul_5_io_vec2_5;
  wire [1:0] VectorMul_5_io_vec2_6;
  wire [1:0] VectorMul_5_io_vec2_7;
  wire [1:0] VectorMul_5_io_vec2_8;
  wire [1:0] VectorMul_5_io_out;
  wire  VectorMul_6_clock;
  wire  VectorMul_6_reset;
  wire [1:0] VectorMul_6_io_vec1_0;
  wire [1:0] VectorMul_6_io_vec1_1;
  wire [1:0] VectorMul_6_io_vec1_2;
  wire [1:0] VectorMul_6_io_vec1_3;
  wire [1:0] VectorMul_6_io_vec1_4;
  wire [1:0] VectorMul_6_io_vec1_5;
  wire [1:0] VectorMul_6_io_vec1_6;
  wire [1:0] VectorMul_6_io_vec1_7;
  wire [1:0] VectorMul_6_io_vec1_8;
  wire [1:0] VectorMul_6_io_vec2_0;
  wire [1:0] VectorMul_6_io_vec2_1;
  wire [1:0] VectorMul_6_io_vec2_2;
  wire [1:0] VectorMul_6_io_vec2_3;
  wire [1:0] VectorMul_6_io_vec2_4;
  wire [1:0] VectorMul_6_io_vec2_5;
  wire [1:0] VectorMul_6_io_vec2_6;
  wire [1:0] VectorMul_6_io_vec2_7;
  wire [1:0] VectorMul_6_io_vec2_8;
  wire [1:0] VectorMul_6_io_out;
  wire  VectorMul_7_clock;
  wire  VectorMul_7_reset;
  wire [1:0] VectorMul_7_io_vec1_0;
  wire [1:0] VectorMul_7_io_vec1_1;
  wire [1:0] VectorMul_7_io_vec1_2;
  wire [1:0] VectorMul_7_io_vec1_3;
  wire [1:0] VectorMul_7_io_vec1_4;
  wire [1:0] VectorMul_7_io_vec1_5;
  wire [1:0] VectorMul_7_io_vec1_6;
  wire [1:0] VectorMul_7_io_vec1_7;
  wire [1:0] VectorMul_7_io_vec1_8;
  wire [1:0] VectorMul_7_io_vec2_0;
  wire [1:0] VectorMul_7_io_vec2_1;
  wire [1:0] VectorMul_7_io_vec2_2;
  wire [1:0] VectorMul_7_io_vec2_3;
  wire [1:0] VectorMul_7_io_vec2_4;
  wire [1:0] VectorMul_7_io_vec2_5;
  wire [1:0] VectorMul_7_io_vec2_6;
  wire [1:0] VectorMul_7_io_vec2_7;
  wire [1:0] VectorMul_7_io_vec2_8;
  wire [1:0] VectorMul_7_io_out;
  wire  VectorMul_8_clock;
  wire  VectorMul_8_reset;
  wire [1:0] VectorMul_8_io_vec1_0;
  wire [1:0] VectorMul_8_io_vec1_1;
  wire [1:0] VectorMul_8_io_vec1_2;
  wire [1:0] VectorMul_8_io_vec1_3;
  wire [1:0] VectorMul_8_io_vec1_4;
  wire [1:0] VectorMul_8_io_vec1_5;
  wire [1:0] VectorMul_8_io_vec1_6;
  wire [1:0] VectorMul_8_io_vec1_7;
  wire [1:0] VectorMul_8_io_vec1_8;
  wire [1:0] VectorMul_8_io_vec2_0;
  wire [1:0] VectorMul_8_io_vec2_1;
  wire [1:0] VectorMul_8_io_vec2_2;
  wire [1:0] VectorMul_8_io_vec2_3;
  wire [1:0] VectorMul_8_io_vec2_4;
  wire [1:0] VectorMul_8_io_vec2_5;
  wire [1:0] VectorMul_8_io_vec2_6;
  wire [1:0] VectorMul_8_io_vec2_7;
  wire [1:0] VectorMul_8_io_vec2_8;
  wire [1:0] VectorMul_8_io_out;
  wire  VectorMul_9_clock;
  wire  VectorMul_9_reset;
  wire [1:0] VectorMul_9_io_vec1_0;
  wire [1:0] VectorMul_9_io_vec1_1;
  wire [1:0] VectorMul_9_io_vec1_2;
  wire [1:0] VectorMul_9_io_vec1_3;
  wire [1:0] VectorMul_9_io_vec1_4;
  wire [1:0] VectorMul_9_io_vec1_5;
  wire [1:0] VectorMul_9_io_vec1_6;
  wire [1:0] VectorMul_9_io_vec1_7;
  wire [1:0] VectorMul_9_io_vec1_8;
  wire [1:0] VectorMul_9_io_vec2_0;
  wire [1:0] VectorMul_9_io_vec2_1;
  wire [1:0] VectorMul_9_io_vec2_2;
  wire [1:0] VectorMul_9_io_vec2_3;
  wire [1:0] VectorMul_9_io_vec2_4;
  wire [1:0] VectorMul_9_io_vec2_5;
  wire [1:0] VectorMul_9_io_vec2_6;
  wire [1:0] VectorMul_9_io_vec2_7;
  wire [1:0] VectorMul_9_io_vec2_8;
  wire [1:0] VectorMul_9_io_out;
  wire  VectorMul_10_clock;
  wire  VectorMul_10_reset;
  wire [1:0] VectorMul_10_io_vec1_0;
  wire [1:0] VectorMul_10_io_vec1_1;
  wire [1:0] VectorMul_10_io_vec1_2;
  wire [1:0] VectorMul_10_io_vec1_3;
  wire [1:0] VectorMul_10_io_vec1_4;
  wire [1:0] VectorMul_10_io_vec1_5;
  wire [1:0] VectorMul_10_io_vec1_6;
  wire [1:0] VectorMul_10_io_vec1_7;
  wire [1:0] VectorMul_10_io_vec1_8;
  wire [1:0] VectorMul_10_io_vec2_0;
  wire [1:0] VectorMul_10_io_vec2_1;
  wire [1:0] VectorMul_10_io_vec2_2;
  wire [1:0] VectorMul_10_io_vec2_3;
  wire [1:0] VectorMul_10_io_vec2_4;
  wire [1:0] VectorMul_10_io_vec2_5;
  wire [1:0] VectorMul_10_io_vec2_6;
  wire [1:0] VectorMul_10_io_vec2_7;
  wire [1:0] VectorMul_10_io_vec2_8;
  wire [1:0] VectorMul_10_io_out;
  wire  VectorMul_11_clock;
  wire  VectorMul_11_reset;
  wire [1:0] VectorMul_11_io_vec1_0;
  wire [1:0] VectorMul_11_io_vec1_1;
  wire [1:0] VectorMul_11_io_vec1_2;
  wire [1:0] VectorMul_11_io_vec1_3;
  wire [1:0] VectorMul_11_io_vec1_4;
  wire [1:0] VectorMul_11_io_vec1_5;
  wire [1:0] VectorMul_11_io_vec1_6;
  wire [1:0] VectorMul_11_io_vec1_7;
  wire [1:0] VectorMul_11_io_vec1_8;
  wire [1:0] VectorMul_11_io_vec2_0;
  wire [1:0] VectorMul_11_io_vec2_1;
  wire [1:0] VectorMul_11_io_vec2_2;
  wire [1:0] VectorMul_11_io_vec2_3;
  wire [1:0] VectorMul_11_io_vec2_4;
  wire [1:0] VectorMul_11_io_vec2_5;
  wire [1:0] VectorMul_11_io_vec2_6;
  wire [1:0] VectorMul_11_io_vec2_7;
  wire [1:0] VectorMul_11_io_vec2_8;
  wire [1:0] VectorMul_11_io_out;
  wire  VectorMul_12_clock;
  wire  VectorMul_12_reset;
  wire [1:0] VectorMul_12_io_vec1_0;
  wire [1:0] VectorMul_12_io_vec1_1;
  wire [1:0] VectorMul_12_io_vec1_2;
  wire [1:0] VectorMul_12_io_vec1_3;
  wire [1:0] VectorMul_12_io_vec1_4;
  wire [1:0] VectorMul_12_io_vec1_5;
  wire [1:0] VectorMul_12_io_vec1_6;
  wire [1:0] VectorMul_12_io_vec1_7;
  wire [1:0] VectorMul_12_io_vec1_8;
  wire [1:0] VectorMul_12_io_vec2_0;
  wire [1:0] VectorMul_12_io_vec2_1;
  wire [1:0] VectorMul_12_io_vec2_2;
  wire [1:0] VectorMul_12_io_vec2_3;
  wire [1:0] VectorMul_12_io_vec2_4;
  wire [1:0] VectorMul_12_io_vec2_5;
  wire [1:0] VectorMul_12_io_vec2_6;
  wire [1:0] VectorMul_12_io_vec2_7;
  wire [1:0] VectorMul_12_io_vec2_8;
  wire [1:0] VectorMul_12_io_out;
  wire  VectorMul_13_clock;
  wire  VectorMul_13_reset;
  wire [1:0] VectorMul_13_io_vec1_0;
  wire [1:0] VectorMul_13_io_vec1_1;
  wire [1:0] VectorMul_13_io_vec1_2;
  wire [1:0] VectorMul_13_io_vec1_3;
  wire [1:0] VectorMul_13_io_vec1_4;
  wire [1:0] VectorMul_13_io_vec1_5;
  wire [1:0] VectorMul_13_io_vec1_6;
  wire [1:0] VectorMul_13_io_vec1_7;
  wire [1:0] VectorMul_13_io_vec1_8;
  wire [1:0] VectorMul_13_io_vec2_0;
  wire [1:0] VectorMul_13_io_vec2_1;
  wire [1:0] VectorMul_13_io_vec2_2;
  wire [1:0] VectorMul_13_io_vec2_3;
  wire [1:0] VectorMul_13_io_vec2_4;
  wire [1:0] VectorMul_13_io_vec2_5;
  wire [1:0] VectorMul_13_io_vec2_6;
  wire [1:0] VectorMul_13_io_vec2_7;
  wire [1:0] VectorMul_13_io_vec2_8;
  wire [1:0] VectorMul_13_io_out;
  wire  VectorMul_14_clock;
  wire  VectorMul_14_reset;
  wire [1:0] VectorMul_14_io_vec1_0;
  wire [1:0] VectorMul_14_io_vec1_1;
  wire [1:0] VectorMul_14_io_vec1_2;
  wire [1:0] VectorMul_14_io_vec1_3;
  wire [1:0] VectorMul_14_io_vec1_4;
  wire [1:0] VectorMul_14_io_vec1_5;
  wire [1:0] VectorMul_14_io_vec1_6;
  wire [1:0] VectorMul_14_io_vec1_7;
  wire [1:0] VectorMul_14_io_vec1_8;
  wire [1:0] VectorMul_14_io_vec2_0;
  wire [1:0] VectorMul_14_io_vec2_1;
  wire [1:0] VectorMul_14_io_vec2_2;
  wire [1:0] VectorMul_14_io_vec2_3;
  wire [1:0] VectorMul_14_io_vec2_4;
  wire [1:0] VectorMul_14_io_vec2_5;
  wire [1:0] VectorMul_14_io_vec2_6;
  wire [1:0] VectorMul_14_io_vec2_7;
  wire [1:0] VectorMul_14_io_vec2_8;
  wire [1:0] VectorMul_14_io_out;
  wire  VectorMul_15_clock;
  wire  VectorMul_15_reset;
  wire [1:0] VectorMul_15_io_vec1_0;
  wire [1:0] VectorMul_15_io_vec1_1;
  wire [1:0] VectorMul_15_io_vec1_2;
  wire [1:0] VectorMul_15_io_vec1_3;
  wire [1:0] VectorMul_15_io_vec1_4;
  wire [1:0] VectorMul_15_io_vec1_5;
  wire [1:0] VectorMul_15_io_vec1_6;
  wire [1:0] VectorMul_15_io_vec1_7;
  wire [1:0] VectorMul_15_io_vec1_8;
  wire [1:0] VectorMul_15_io_vec2_0;
  wire [1:0] VectorMul_15_io_vec2_1;
  wire [1:0] VectorMul_15_io_vec2_2;
  wire [1:0] VectorMul_15_io_vec2_3;
  wire [1:0] VectorMul_15_io_vec2_4;
  wire [1:0] VectorMul_15_io_vec2_5;
  wire [1:0] VectorMul_15_io_vec2_6;
  wire [1:0] VectorMul_15_io_vec2_7;
  wire [1:0] VectorMul_15_io_vec2_8;
  wire [1:0] VectorMul_15_io_out;
  wire  VectorMul_16_clock;
  wire  VectorMul_16_reset;
  wire [1:0] VectorMul_16_io_vec1_0;
  wire [1:0] VectorMul_16_io_vec1_1;
  wire [1:0] VectorMul_16_io_vec1_2;
  wire [1:0] VectorMul_16_io_vec1_3;
  wire [1:0] VectorMul_16_io_vec1_4;
  wire [1:0] VectorMul_16_io_vec1_5;
  wire [1:0] VectorMul_16_io_vec1_6;
  wire [1:0] VectorMul_16_io_vec1_7;
  wire [1:0] VectorMul_16_io_vec1_8;
  wire [1:0] VectorMul_16_io_vec2_0;
  wire [1:0] VectorMul_16_io_vec2_1;
  wire [1:0] VectorMul_16_io_vec2_2;
  wire [1:0] VectorMul_16_io_vec2_3;
  wire [1:0] VectorMul_16_io_vec2_4;
  wire [1:0] VectorMul_16_io_vec2_5;
  wire [1:0] VectorMul_16_io_vec2_6;
  wire [1:0] VectorMul_16_io_vec2_7;
  wire [1:0] VectorMul_16_io_vec2_8;
  wire [1:0] VectorMul_16_io_out;
  wire  VectorMul_17_clock;
  wire  VectorMul_17_reset;
  wire [1:0] VectorMul_17_io_vec1_0;
  wire [1:0] VectorMul_17_io_vec1_1;
  wire [1:0] VectorMul_17_io_vec1_2;
  wire [1:0] VectorMul_17_io_vec1_3;
  wire [1:0] VectorMul_17_io_vec1_4;
  wire [1:0] VectorMul_17_io_vec1_5;
  wire [1:0] VectorMul_17_io_vec1_6;
  wire [1:0] VectorMul_17_io_vec1_7;
  wire [1:0] VectorMul_17_io_vec1_8;
  wire [1:0] VectorMul_17_io_vec2_0;
  wire [1:0] VectorMul_17_io_vec2_1;
  wire [1:0] VectorMul_17_io_vec2_2;
  wire [1:0] VectorMul_17_io_vec2_3;
  wire [1:0] VectorMul_17_io_vec2_4;
  wire [1:0] VectorMul_17_io_vec2_5;
  wire [1:0] VectorMul_17_io_vec2_6;
  wire [1:0] VectorMul_17_io_vec2_7;
  wire [1:0] VectorMul_17_io_vec2_8;
  wire [1:0] VectorMul_17_io_out;
  wire  VectorMul_18_clock;
  wire  VectorMul_18_reset;
  wire [1:0] VectorMul_18_io_vec1_0;
  wire [1:0] VectorMul_18_io_vec1_1;
  wire [1:0] VectorMul_18_io_vec1_2;
  wire [1:0] VectorMul_18_io_vec1_3;
  wire [1:0] VectorMul_18_io_vec1_4;
  wire [1:0] VectorMul_18_io_vec1_5;
  wire [1:0] VectorMul_18_io_vec1_6;
  wire [1:0] VectorMul_18_io_vec1_7;
  wire [1:0] VectorMul_18_io_vec1_8;
  wire [1:0] VectorMul_18_io_vec2_0;
  wire [1:0] VectorMul_18_io_vec2_1;
  wire [1:0] VectorMul_18_io_vec2_2;
  wire [1:0] VectorMul_18_io_vec2_3;
  wire [1:0] VectorMul_18_io_vec2_4;
  wire [1:0] VectorMul_18_io_vec2_5;
  wire [1:0] VectorMul_18_io_vec2_6;
  wire [1:0] VectorMul_18_io_vec2_7;
  wire [1:0] VectorMul_18_io_vec2_8;
  wire [1:0] VectorMul_18_io_out;
  wire  VectorMul_19_clock;
  wire  VectorMul_19_reset;
  wire [1:0] VectorMul_19_io_vec1_0;
  wire [1:0] VectorMul_19_io_vec1_1;
  wire [1:0] VectorMul_19_io_vec1_2;
  wire [1:0] VectorMul_19_io_vec1_3;
  wire [1:0] VectorMul_19_io_vec1_4;
  wire [1:0] VectorMul_19_io_vec1_5;
  wire [1:0] VectorMul_19_io_vec1_6;
  wire [1:0] VectorMul_19_io_vec1_7;
  wire [1:0] VectorMul_19_io_vec1_8;
  wire [1:0] VectorMul_19_io_vec2_0;
  wire [1:0] VectorMul_19_io_vec2_1;
  wire [1:0] VectorMul_19_io_vec2_2;
  wire [1:0] VectorMul_19_io_vec2_3;
  wire [1:0] VectorMul_19_io_vec2_4;
  wire [1:0] VectorMul_19_io_vec2_5;
  wire [1:0] VectorMul_19_io_vec2_6;
  wire [1:0] VectorMul_19_io_vec2_7;
  wire [1:0] VectorMul_19_io_vec2_8;
  wire [1:0] VectorMul_19_io_out;
  wire  VectorMul_20_clock;
  wire  VectorMul_20_reset;
  wire [1:0] VectorMul_20_io_vec1_0;
  wire [1:0] VectorMul_20_io_vec1_1;
  wire [1:0] VectorMul_20_io_vec1_2;
  wire [1:0] VectorMul_20_io_vec1_3;
  wire [1:0] VectorMul_20_io_vec1_4;
  wire [1:0] VectorMul_20_io_vec1_5;
  wire [1:0] VectorMul_20_io_vec1_6;
  wire [1:0] VectorMul_20_io_vec1_7;
  wire [1:0] VectorMul_20_io_vec1_8;
  wire [1:0] VectorMul_20_io_vec2_0;
  wire [1:0] VectorMul_20_io_vec2_1;
  wire [1:0] VectorMul_20_io_vec2_2;
  wire [1:0] VectorMul_20_io_vec2_3;
  wire [1:0] VectorMul_20_io_vec2_4;
  wire [1:0] VectorMul_20_io_vec2_5;
  wire [1:0] VectorMul_20_io_vec2_6;
  wire [1:0] VectorMul_20_io_vec2_7;
  wire [1:0] VectorMul_20_io_vec2_8;
  wire [1:0] VectorMul_20_io_out;
  wire  VectorMul_21_clock;
  wire  VectorMul_21_reset;
  wire [1:0] VectorMul_21_io_vec1_0;
  wire [1:0] VectorMul_21_io_vec1_1;
  wire [1:0] VectorMul_21_io_vec1_2;
  wire [1:0] VectorMul_21_io_vec1_3;
  wire [1:0] VectorMul_21_io_vec1_4;
  wire [1:0] VectorMul_21_io_vec1_5;
  wire [1:0] VectorMul_21_io_vec1_6;
  wire [1:0] VectorMul_21_io_vec1_7;
  wire [1:0] VectorMul_21_io_vec1_8;
  wire [1:0] VectorMul_21_io_vec2_0;
  wire [1:0] VectorMul_21_io_vec2_1;
  wire [1:0] VectorMul_21_io_vec2_2;
  wire [1:0] VectorMul_21_io_vec2_3;
  wire [1:0] VectorMul_21_io_vec2_4;
  wire [1:0] VectorMul_21_io_vec2_5;
  wire [1:0] VectorMul_21_io_vec2_6;
  wire [1:0] VectorMul_21_io_vec2_7;
  wire [1:0] VectorMul_21_io_vec2_8;
  wire [1:0] VectorMul_21_io_out;
  wire  VectorMul_22_clock;
  wire  VectorMul_22_reset;
  wire [1:0] VectorMul_22_io_vec1_0;
  wire [1:0] VectorMul_22_io_vec1_1;
  wire [1:0] VectorMul_22_io_vec1_2;
  wire [1:0] VectorMul_22_io_vec1_3;
  wire [1:0] VectorMul_22_io_vec1_4;
  wire [1:0] VectorMul_22_io_vec1_5;
  wire [1:0] VectorMul_22_io_vec1_6;
  wire [1:0] VectorMul_22_io_vec1_7;
  wire [1:0] VectorMul_22_io_vec1_8;
  wire [1:0] VectorMul_22_io_vec2_0;
  wire [1:0] VectorMul_22_io_vec2_1;
  wire [1:0] VectorMul_22_io_vec2_2;
  wire [1:0] VectorMul_22_io_vec2_3;
  wire [1:0] VectorMul_22_io_vec2_4;
  wire [1:0] VectorMul_22_io_vec2_5;
  wire [1:0] VectorMul_22_io_vec2_6;
  wire [1:0] VectorMul_22_io_vec2_7;
  wire [1:0] VectorMul_22_io_vec2_8;
  wire [1:0] VectorMul_22_io_out;
  wire  VectorMul_23_clock;
  wire  VectorMul_23_reset;
  wire [1:0] VectorMul_23_io_vec1_0;
  wire [1:0] VectorMul_23_io_vec1_1;
  wire [1:0] VectorMul_23_io_vec1_2;
  wire [1:0] VectorMul_23_io_vec1_3;
  wire [1:0] VectorMul_23_io_vec1_4;
  wire [1:0] VectorMul_23_io_vec1_5;
  wire [1:0] VectorMul_23_io_vec1_6;
  wire [1:0] VectorMul_23_io_vec1_7;
  wire [1:0] VectorMul_23_io_vec1_8;
  wire [1:0] VectorMul_23_io_vec2_0;
  wire [1:0] VectorMul_23_io_vec2_1;
  wire [1:0] VectorMul_23_io_vec2_2;
  wire [1:0] VectorMul_23_io_vec2_3;
  wire [1:0] VectorMul_23_io_vec2_4;
  wire [1:0] VectorMul_23_io_vec2_5;
  wire [1:0] VectorMul_23_io_vec2_6;
  wire [1:0] VectorMul_23_io_vec2_7;
  wire [1:0] VectorMul_23_io_vec2_8;
  wire [1:0] VectorMul_23_io_out;
  wire  VectorMul_24_clock;
  wire  VectorMul_24_reset;
  wire [1:0] VectorMul_24_io_vec1_0;
  wire [1:0] VectorMul_24_io_vec1_1;
  wire [1:0] VectorMul_24_io_vec1_2;
  wire [1:0] VectorMul_24_io_vec1_3;
  wire [1:0] VectorMul_24_io_vec1_4;
  wire [1:0] VectorMul_24_io_vec1_5;
  wire [1:0] VectorMul_24_io_vec1_6;
  wire [1:0] VectorMul_24_io_vec1_7;
  wire [1:0] VectorMul_24_io_vec1_8;
  wire [1:0] VectorMul_24_io_vec2_0;
  wire [1:0] VectorMul_24_io_vec2_1;
  wire [1:0] VectorMul_24_io_vec2_2;
  wire [1:0] VectorMul_24_io_vec2_3;
  wire [1:0] VectorMul_24_io_vec2_4;
  wire [1:0] VectorMul_24_io_vec2_5;
  wire [1:0] VectorMul_24_io_vec2_6;
  wire [1:0] VectorMul_24_io_vec2_7;
  wire [1:0] VectorMul_24_io_vec2_8;
  wire [1:0] VectorMul_24_io_out;
  wire [1:0] result_0;
  wire [1:0] result_1;
  wire [1:0] result_2;
  wire [1:0] result_3;
  wire [1:0] result_4;
  wire [1:0] result_5;
  wire [1:0] result_6;
  wire [1:0] result_7;
  wire [1:0] result_8;
  wire [1:0] result_9;
  wire [1:0] result_10;
  wire [1:0] result_11;
  wire [1:0] result_12;
  wire [1:0] result_13;
  wire [1:0] result_14;
  wire [1:0] result_15;
  wire [1:0] result_16;
  wire [1:0] result_17;
  wire [1:0] result_18;
  wire [1:0] result_19;
  wire [1:0] result_20;
  wire [1:0] result_21;
  wire [1:0] result_22;
  wire [1:0] result_23;
  wire [1:0] result_24;
  reg [1:0] xx_8;
  reg [31:0] _RAND_0;
  reg [1:0] xx_9;
  reg [31:0] _RAND_1;
  reg [1:0] xx_10;
  reg [31:0] _RAND_2;
  reg [1:0] xx_11;
  reg [31:0] _RAND_3;
  reg [1:0] xx_12;
  reg [31:0] _RAND_4;
  reg [1:0] xx_15;
  reg [31:0] _RAND_5;
  reg [1:0] xx_16;
  reg [31:0] _RAND_6;
  reg [1:0] xx_17;
  reg [31:0] _RAND_7;
  reg [1:0] xx_18;
  reg [31:0] _RAND_8;
  reg [1:0] xx_19;
  reg [31:0] _RAND_9;
  reg [1:0] xx_22;
  reg [31:0] _RAND_10;
  reg [1:0] xx_23;
  reg [31:0] _RAND_11;
  reg [1:0] xx_24;
  reg [31:0] _RAND_12;
  reg [1:0] xx_25;
  reg [31:0] _RAND_13;
  reg [1:0] xx_26;
  reg [31:0] _RAND_14;
  reg [1:0] xx_29;
  reg [31:0] _RAND_15;
  reg [1:0] xx_30;
  reg [31:0] _RAND_16;
  reg [1:0] xx_31;
  reg [31:0] _RAND_17;
  reg [1:0] xx_32;
  reg [31:0] _RAND_18;
  reg [1:0] xx_33;
  reg [31:0] _RAND_19;
  reg [1:0] xx_36;
  reg [31:0] _RAND_20;
  reg [1:0] xx_37;
  reg [31:0] _RAND_21;
  reg [1:0] xx_38;
  reg [31:0] _RAND_22;
  reg [1:0] xx_39;
  reg [31:0] _RAND_23;
  reg [1:0] xx_40;
  reg [31:0] _RAND_24;
  reg [1:0] _T_507_4;
  reg [31:0] _RAND_25;
  reg [1:0] _T_507_5;
  reg [31:0] _RAND_26;
  reg [1:0] _T_507_7;
  reg [31:0] _RAND_27;
  reg [1:0] _T_507_8;
  reg [31:0] _RAND_28;
  reg [1:0] _T_584_1;
  reg [31:0] _RAND_29;
  reg [1:0] _T_584_2;
  reg [31:0] _RAND_30;
  reg [1:0] _T_584_4;
  reg [31:0] _RAND_31;
  reg [1:0] _T_584_5;
  reg [31:0] _RAND_32;
  reg [1:0] _T_584_7;
  reg [31:0] _RAND_33;
  reg [1:0] _T_584_8;
  reg [31:0] _RAND_34;
  reg [1:0] _T_661_1;
  reg [31:0] _RAND_35;
  reg [1:0] _T_661_2;
  reg [31:0] _RAND_36;
  reg [1:0] _T_661_4;
  reg [31:0] _RAND_37;
  reg [1:0] _T_661_5;
  reg [31:0] _RAND_38;
  reg [1:0] _T_661_7;
  reg [31:0] _RAND_39;
  reg [1:0] _T_661_8;
  reg [31:0] _RAND_40;
  reg [1:0] _T_738_1;
  reg [31:0] _RAND_41;
  reg [1:0] _T_738_2;
  reg [31:0] _RAND_42;
  reg [1:0] _T_738_4;
  reg [31:0] _RAND_43;
  reg [1:0] _T_738_5;
  reg [31:0] _RAND_44;
  reg [1:0] _T_738_7;
  reg [31:0] _RAND_45;
  reg [1:0] _T_738_8;
  reg [31:0] _RAND_46;
  reg [1:0] _T_815_1;
  reg [31:0] _RAND_47;
  reg [1:0] _T_815_2;
  reg [31:0] _RAND_48;
  reg [1:0] _T_815_4;
  reg [31:0] _RAND_49;
  reg [1:0] _T_815_5;
  reg [31:0] _RAND_50;
  reg [1:0] _T_892_3;
  reg [31:0] _RAND_51;
  reg [1:0] _T_892_4;
  reg [31:0] _RAND_52;
  reg [1:0] _T_892_5;
  reg [31:0] _RAND_53;
  reg [1:0] _T_892_6;
  reg [31:0] _RAND_54;
  reg [1:0] _T_892_7;
  reg [31:0] _RAND_55;
  reg [1:0] _T_892_8;
  reg [31:0] _RAND_56;
  reg [1:0] _T_969_0;
  reg [31:0] _RAND_57;
  reg [1:0] _T_969_1;
  reg [31:0] _RAND_58;
  reg [1:0] _T_969_2;
  reg [31:0] _RAND_59;
  reg [1:0] _T_969_3;
  reg [31:0] _RAND_60;
  reg [1:0] _T_969_4;
  reg [31:0] _RAND_61;
  reg [1:0] _T_969_5;
  reg [31:0] _RAND_62;
  reg [1:0] _T_969_6;
  reg [31:0] _RAND_63;
  reg [1:0] _T_969_7;
  reg [31:0] _RAND_64;
  reg [1:0] _T_969_8;
  reg [31:0] _RAND_65;
  reg [1:0] _T_1046_0;
  reg [31:0] _RAND_66;
  reg [1:0] _T_1046_1;
  reg [31:0] _RAND_67;
  reg [1:0] _T_1046_2;
  reg [31:0] _RAND_68;
  reg [1:0] _T_1046_3;
  reg [31:0] _RAND_69;
  reg [1:0] _T_1046_4;
  reg [31:0] _RAND_70;
  reg [1:0] _T_1046_5;
  reg [31:0] _RAND_71;
  reg [1:0] _T_1046_6;
  reg [31:0] _RAND_72;
  reg [1:0] _T_1046_7;
  reg [31:0] _RAND_73;
  reg [1:0] _T_1046_8;
  reg [31:0] _RAND_74;
  reg [1:0] _T_1123_0;
  reg [31:0] _RAND_75;
  reg [1:0] _T_1123_1;
  reg [31:0] _RAND_76;
  reg [1:0] _T_1123_2;
  reg [31:0] _RAND_77;
  reg [1:0] _T_1123_3;
  reg [31:0] _RAND_78;
  reg [1:0] _T_1123_4;
  reg [31:0] _RAND_79;
  reg [1:0] _T_1123_5;
  reg [31:0] _RAND_80;
  reg [1:0] _T_1123_6;
  reg [31:0] _RAND_81;
  reg [1:0] _T_1123_7;
  reg [31:0] _RAND_82;
  reg [1:0] _T_1123_8;
  reg [31:0] _RAND_83;
  reg [1:0] _T_1200_0;
  reg [31:0] _RAND_84;
  reg [1:0] _T_1200_1;
  reg [31:0] _RAND_85;
  reg [1:0] _T_1200_2;
  reg [31:0] _RAND_86;
  reg [1:0] _T_1200_3;
  reg [31:0] _RAND_87;
  reg [1:0] _T_1200_4;
  reg [31:0] _RAND_88;
  reg [1:0] _T_1200_5;
  reg [31:0] _RAND_89;
  reg [1:0] _T_1277_3;
  reg [31:0] _RAND_90;
  reg [1:0] _T_1277_4;
  reg [31:0] _RAND_91;
  reg [1:0] _T_1277_5;
  reg [31:0] _RAND_92;
  reg [1:0] _T_1277_6;
  reg [31:0] _RAND_93;
  reg [1:0] _T_1277_7;
  reg [31:0] _RAND_94;
  reg [1:0] _T_1277_8;
  reg [31:0] _RAND_95;
  reg [1:0] _T_1354_0;
  reg [31:0] _RAND_96;
  reg [1:0] _T_1354_1;
  reg [31:0] _RAND_97;
  reg [1:0] _T_1354_2;
  reg [31:0] _RAND_98;
  reg [1:0] _T_1354_3;
  reg [31:0] _RAND_99;
  reg [1:0] _T_1354_4;
  reg [31:0] _RAND_100;
  reg [1:0] _T_1354_5;
  reg [31:0] _RAND_101;
  reg [1:0] _T_1354_6;
  reg [31:0] _RAND_102;
  reg [1:0] _T_1354_7;
  reg [31:0] _RAND_103;
  reg [1:0] _T_1354_8;
  reg [31:0] _RAND_104;
  reg [1:0] _T_1431_0;
  reg [31:0] _RAND_105;
  reg [1:0] _T_1431_1;
  reg [31:0] _RAND_106;
  reg [1:0] _T_1431_2;
  reg [31:0] _RAND_107;
  reg [1:0] _T_1431_3;
  reg [31:0] _RAND_108;
  reg [1:0] _T_1431_4;
  reg [31:0] _RAND_109;
  reg [1:0] _T_1431_5;
  reg [31:0] _RAND_110;
  reg [1:0] _T_1431_6;
  reg [31:0] _RAND_111;
  reg [1:0] _T_1431_7;
  reg [31:0] _RAND_112;
  reg [1:0] _T_1431_8;
  reg [31:0] _RAND_113;
  reg [1:0] _T_1508_0;
  reg [31:0] _RAND_114;
  reg [1:0] _T_1508_1;
  reg [31:0] _RAND_115;
  reg [1:0] _T_1508_2;
  reg [31:0] _RAND_116;
  reg [1:0] _T_1508_3;
  reg [31:0] _RAND_117;
  reg [1:0] _T_1508_4;
  reg [31:0] _RAND_118;
  reg [1:0] _T_1508_5;
  reg [31:0] _RAND_119;
  reg [1:0] _T_1508_6;
  reg [31:0] _RAND_120;
  reg [1:0] _T_1508_7;
  reg [31:0] _RAND_121;
  reg [1:0] _T_1508_8;
  reg [31:0] _RAND_122;
  reg [1:0] _T_1585_0;
  reg [31:0] _RAND_123;
  reg [1:0] _T_1585_1;
  reg [31:0] _RAND_124;
  reg [1:0] _T_1585_2;
  reg [31:0] _RAND_125;
  reg [1:0] _T_1585_3;
  reg [31:0] _RAND_126;
  reg [1:0] _T_1585_4;
  reg [31:0] _RAND_127;
  reg [1:0] _T_1585_5;
  reg [31:0] _RAND_128;
  reg [1:0] _T_1662_3;
  reg [31:0] _RAND_129;
  reg [1:0] _T_1662_4;
  reg [31:0] _RAND_130;
  reg [1:0] _T_1662_5;
  reg [31:0] _RAND_131;
  reg [1:0] _T_1662_6;
  reg [31:0] _RAND_132;
  reg [1:0] _T_1662_7;
  reg [31:0] _RAND_133;
  reg [1:0] _T_1662_8;
  reg [31:0] _RAND_134;
  reg [1:0] _T_1739_0;
  reg [31:0] _RAND_135;
  reg [1:0] _T_1739_1;
  reg [31:0] _RAND_136;
  reg [1:0] _T_1739_2;
  reg [31:0] _RAND_137;
  reg [1:0] _T_1739_3;
  reg [31:0] _RAND_138;
  reg [1:0] _T_1739_4;
  reg [31:0] _RAND_139;
  reg [1:0] _T_1739_5;
  reg [31:0] _RAND_140;
  reg [1:0] _T_1739_6;
  reg [31:0] _RAND_141;
  reg [1:0] _T_1739_7;
  reg [31:0] _RAND_142;
  reg [1:0] _T_1739_8;
  reg [31:0] _RAND_143;
  reg [1:0] _T_1816_0;
  reg [31:0] _RAND_144;
  reg [1:0] _T_1816_1;
  reg [31:0] _RAND_145;
  reg [1:0] _T_1816_2;
  reg [31:0] _RAND_146;
  reg [1:0] _T_1816_3;
  reg [31:0] _RAND_147;
  reg [1:0] _T_1816_4;
  reg [31:0] _RAND_148;
  reg [1:0] _T_1816_5;
  reg [31:0] _RAND_149;
  reg [1:0] _T_1816_6;
  reg [31:0] _RAND_150;
  reg [1:0] _T_1816_7;
  reg [31:0] _RAND_151;
  reg [1:0] _T_1816_8;
  reg [31:0] _RAND_152;
  reg [1:0] _T_1893_0;
  reg [31:0] _RAND_153;
  reg [1:0] _T_1893_1;
  reg [31:0] _RAND_154;
  reg [1:0] _T_1893_2;
  reg [31:0] _RAND_155;
  reg [1:0] _T_1893_3;
  reg [31:0] _RAND_156;
  reg [1:0] _T_1893_4;
  reg [31:0] _RAND_157;
  reg [1:0] _T_1893_5;
  reg [31:0] _RAND_158;
  reg [1:0] _T_1893_6;
  reg [31:0] _RAND_159;
  reg [1:0] _T_1893_7;
  reg [31:0] _RAND_160;
  reg [1:0] _T_1893_8;
  reg [31:0] _RAND_161;
  reg [1:0] _T_1970_0;
  reg [31:0] _RAND_162;
  reg [1:0] _T_1970_1;
  reg [31:0] _RAND_163;
  reg [1:0] _T_1970_2;
  reg [31:0] _RAND_164;
  reg [1:0] _T_1970_3;
  reg [31:0] _RAND_165;
  reg [1:0] _T_1970_4;
  reg [31:0] _RAND_166;
  reg [1:0] _T_1970_5;
  reg [31:0] _RAND_167;
  reg [1:0] _T_2047_3;
  reg [31:0] _RAND_168;
  reg [1:0] _T_2047_4;
  reg [31:0] _RAND_169;
  reg [1:0] _T_2047_6;
  reg [31:0] _RAND_170;
  reg [1:0] _T_2047_7;
  reg [31:0] _RAND_171;
  reg [1:0] _T_2124_0;
  reg [31:0] _RAND_172;
  reg [1:0] _T_2124_1;
  reg [31:0] _RAND_173;
  reg [1:0] _T_2124_3;
  reg [31:0] _RAND_174;
  reg [1:0] _T_2124_4;
  reg [31:0] _RAND_175;
  reg [1:0] _T_2124_6;
  reg [31:0] _RAND_176;
  reg [1:0] _T_2124_7;
  reg [31:0] _RAND_177;
  reg [1:0] _T_2201_0;
  reg [31:0] _RAND_178;
  reg [1:0] _T_2201_1;
  reg [31:0] _RAND_179;
  reg [1:0] _T_2201_3;
  reg [31:0] _RAND_180;
  reg [1:0] _T_2201_4;
  reg [31:0] _RAND_181;
  reg [1:0] _T_2201_6;
  reg [31:0] _RAND_182;
  reg [1:0] _T_2201_7;
  reg [31:0] _RAND_183;
  reg [1:0] _T_2278_0;
  reg [31:0] _RAND_184;
  reg [1:0] _T_2278_1;
  reg [31:0] _RAND_185;
  reg [1:0] _T_2278_3;
  reg [31:0] _RAND_186;
  reg [1:0] _T_2278_4;
  reg [31:0] _RAND_187;
  reg [1:0] _T_2278_6;
  reg [31:0] _RAND_188;
  reg [1:0] _T_2278_7;
  reg [31:0] _RAND_189;
  reg [1:0] _T_2355_0;
  reg [31:0] _RAND_190;
  reg [1:0] _T_2355_1;
  reg [31:0] _RAND_191;
  reg [1:0] _T_2355_3;
  reg [31:0] _RAND_192;
  reg [1:0] _T_2355_4;
  reg [31:0] _RAND_193;
  VectorMul VectorMul (
    .clock(VectorMul_clock),
    .reset(VectorMul_reset),
    .io_vec1_0(VectorMul_io_vec1_0),
    .io_vec1_1(VectorMul_io_vec1_1),
    .io_vec1_2(VectorMul_io_vec1_2),
    .io_vec1_3(VectorMul_io_vec1_3),
    .io_vec1_4(VectorMul_io_vec1_4),
    .io_vec1_5(VectorMul_io_vec1_5),
    .io_vec1_6(VectorMul_io_vec1_6),
    .io_vec1_7(VectorMul_io_vec1_7),
    .io_vec1_8(VectorMul_io_vec1_8),
    .io_vec2_0(VectorMul_io_vec2_0),
    .io_vec2_1(VectorMul_io_vec2_1),
    .io_vec2_2(VectorMul_io_vec2_2),
    .io_vec2_3(VectorMul_io_vec2_3),
    .io_vec2_4(VectorMul_io_vec2_4),
    .io_vec2_5(VectorMul_io_vec2_5),
    .io_vec2_6(VectorMul_io_vec2_6),
    .io_vec2_7(VectorMul_io_vec2_7),
    .io_vec2_8(VectorMul_io_vec2_8),
    .io_out(VectorMul_io_out)
  );
  VectorMul VectorMul_1 (
    .clock(VectorMul_1_clock),
    .reset(VectorMul_1_reset),
    .io_vec1_0(VectorMul_1_io_vec1_0),
    .io_vec1_1(VectorMul_1_io_vec1_1),
    .io_vec1_2(VectorMul_1_io_vec1_2),
    .io_vec1_3(VectorMul_1_io_vec1_3),
    .io_vec1_4(VectorMul_1_io_vec1_4),
    .io_vec1_5(VectorMul_1_io_vec1_5),
    .io_vec1_6(VectorMul_1_io_vec1_6),
    .io_vec1_7(VectorMul_1_io_vec1_7),
    .io_vec1_8(VectorMul_1_io_vec1_8),
    .io_vec2_0(VectorMul_1_io_vec2_0),
    .io_vec2_1(VectorMul_1_io_vec2_1),
    .io_vec2_2(VectorMul_1_io_vec2_2),
    .io_vec2_3(VectorMul_1_io_vec2_3),
    .io_vec2_4(VectorMul_1_io_vec2_4),
    .io_vec2_5(VectorMul_1_io_vec2_5),
    .io_vec2_6(VectorMul_1_io_vec2_6),
    .io_vec2_7(VectorMul_1_io_vec2_7),
    .io_vec2_8(VectorMul_1_io_vec2_8),
    .io_out(VectorMul_1_io_out)
  );
  VectorMul VectorMul_2 (
    .clock(VectorMul_2_clock),
    .reset(VectorMul_2_reset),
    .io_vec1_0(VectorMul_2_io_vec1_0),
    .io_vec1_1(VectorMul_2_io_vec1_1),
    .io_vec1_2(VectorMul_2_io_vec1_2),
    .io_vec1_3(VectorMul_2_io_vec1_3),
    .io_vec1_4(VectorMul_2_io_vec1_4),
    .io_vec1_5(VectorMul_2_io_vec1_5),
    .io_vec1_6(VectorMul_2_io_vec1_6),
    .io_vec1_7(VectorMul_2_io_vec1_7),
    .io_vec1_8(VectorMul_2_io_vec1_8),
    .io_vec2_0(VectorMul_2_io_vec2_0),
    .io_vec2_1(VectorMul_2_io_vec2_1),
    .io_vec2_2(VectorMul_2_io_vec2_2),
    .io_vec2_3(VectorMul_2_io_vec2_3),
    .io_vec2_4(VectorMul_2_io_vec2_4),
    .io_vec2_5(VectorMul_2_io_vec2_5),
    .io_vec2_6(VectorMul_2_io_vec2_6),
    .io_vec2_7(VectorMul_2_io_vec2_7),
    .io_vec2_8(VectorMul_2_io_vec2_8),
    .io_out(VectorMul_2_io_out)
  );
  VectorMul VectorMul_3 (
    .clock(VectorMul_3_clock),
    .reset(VectorMul_3_reset),
    .io_vec1_0(VectorMul_3_io_vec1_0),
    .io_vec1_1(VectorMul_3_io_vec1_1),
    .io_vec1_2(VectorMul_3_io_vec1_2),
    .io_vec1_3(VectorMul_3_io_vec1_3),
    .io_vec1_4(VectorMul_3_io_vec1_4),
    .io_vec1_5(VectorMul_3_io_vec1_5),
    .io_vec1_6(VectorMul_3_io_vec1_6),
    .io_vec1_7(VectorMul_3_io_vec1_7),
    .io_vec1_8(VectorMul_3_io_vec1_8),
    .io_vec2_0(VectorMul_3_io_vec2_0),
    .io_vec2_1(VectorMul_3_io_vec2_1),
    .io_vec2_2(VectorMul_3_io_vec2_2),
    .io_vec2_3(VectorMul_3_io_vec2_3),
    .io_vec2_4(VectorMul_3_io_vec2_4),
    .io_vec2_5(VectorMul_3_io_vec2_5),
    .io_vec2_6(VectorMul_3_io_vec2_6),
    .io_vec2_7(VectorMul_3_io_vec2_7),
    .io_vec2_8(VectorMul_3_io_vec2_8),
    .io_out(VectorMul_3_io_out)
  );
  VectorMul VectorMul_4 (
    .clock(VectorMul_4_clock),
    .reset(VectorMul_4_reset),
    .io_vec1_0(VectorMul_4_io_vec1_0),
    .io_vec1_1(VectorMul_4_io_vec1_1),
    .io_vec1_2(VectorMul_4_io_vec1_2),
    .io_vec1_3(VectorMul_4_io_vec1_3),
    .io_vec1_4(VectorMul_4_io_vec1_4),
    .io_vec1_5(VectorMul_4_io_vec1_5),
    .io_vec1_6(VectorMul_4_io_vec1_6),
    .io_vec1_7(VectorMul_4_io_vec1_7),
    .io_vec1_8(VectorMul_4_io_vec1_8),
    .io_vec2_0(VectorMul_4_io_vec2_0),
    .io_vec2_1(VectorMul_4_io_vec2_1),
    .io_vec2_2(VectorMul_4_io_vec2_2),
    .io_vec2_3(VectorMul_4_io_vec2_3),
    .io_vec2_4(VectorMul_4_io_vec2_4),
    .io_vec2_5(VectorMul_4_io_vec2_5),
    .io_vec2_6(VectorMul_4_io_vec2_6),
    .io_vec2_7(VectorMul_4_io_vec2_7),
    .io_vec2_8(VectorMul_4_io_vec2_8),
    .io_out(VectorMul_4_io_out)
  );
  VectorMul VectorMul_5 (
    .clock(VectorMul_5_clock),
    .reset(VectorMul_5_reset),
    .io_vec1_0(VectorMul_5_io_vec1_0),
    .io_vec1_1(VectorMul_5_io_vec1_1),
    .io_vec1_2(VectorMul_5_io_vec1_2),
    .io_vec1_3(VectorMul_5_io_vec1_3),
    .io_vec1_4(VectorMul_5_io_vec1_4),
    .io_vec1_5(VectorMul_5_io_vec1_5),
    .io_vec1_6(VectorMul_5_io_vec1_6),
    .io_vec1_7(VectorMul_5_io_vec1_7),
    .io_vec1_8(VectorMul_5_io_vec1_8),
    .io_vec2_0(VectorMul_5_io_vec2_0),
    .io_vec2_1(VectorMul_5_io_vec2_1),
    .io_vec2_2(VectorMul_5_io_vec2_2),
    .io_vec2_3(VectorMul_5_io_vec2_3),
    .io_vec2_4(VectorMul_5_io_vec2_4),
    .io_vec2_5(VectorMul_5_io_vec2_5),
    .io_vec2_6(VectorMul_5_io_vec2_6),
    .io_vec2_7(VectorMul_5_io_vec2_7),
    .io_vec2_8(VectorMul_5_io_vec2_8),
    .io_out(VectorMul_5_io_out)
  );
  VectorMul VectorMul_6 (
    .clock(VectorMul_6_clock),
    .reset(VectorMul_6_reset),
    .io_vec1_0(VectorMul_6_io_vec1_0),
    .io_vec1_1(VectorMul_6_io_vec1_1),
    .io_vec1_2(VectorMul_6_io_vec1_2),
    .io_vec1_3(VectorMul_6_io_vec1_3),
    .io_vec1_4(VectorMul_6_io_vec1_4),
    .io_vec1_5(VectorMul_6_io_vec1_5),
    .io_vec1_6(VectorMul_6_io_vec1_6),
    .io_vec1_7(VectorMul_6_io_vec1_7),
    .io_vec1_8(VectorMul_6_io_vec1_8),
    .io_vec2_0(VectorMul_6_io_vec2_0),
    .io_vec2_1(VectorMul_6_io_vec2_1),
    .io_vec2_2(VectorMul_6_io_vec2_2),
    .io_vec2_3(VectorMul_6_io_vec2_3),
    .io_vec2_4(VectorMul_6_io_vec2_4),
    .io_vec2_5(VectorMul_6_io_vec2_5),
    .io_vec2_6(VectorMul_6_io_vec2_6),
    .io_vec2_7(VectorMul_6_io_vec2_7),
    .io_vec2_8(VectorMul_6_io_vec2_8),
    .io_out(VectorMul_6_io_out)
  );
  VectorMul VectorMul_7 (
    .clock(VectorMul_7_clock),
    .reset(VectorMul_7_reset),
    .io_vec1_0(VectorMul_7_io_vec1_0),
    .io_vec1_1(VectorMul_7_io_vec1_1),
    .io_vec1_2(VectorMul_7_io_vec1_2),
    .io_vec1_3(VectorMul_7_io_vec1_3),
    .io_vec1_4(VectorMul_7_io_vec1_4),
    .io_vec1_5(VectorMul_7_io_vec1_5),
    .io_vec1_6(VectorMul_7_io_vec1_6),
    .io_vec1_7(VectorMul_7_io_vec1_7),
    .io_vec1_8(VectorMul_7_io_vec1_8),
    .io_vec2_0(VectorMul_7_io_vec2_0),
    .io_vec2_1(VectorMul_7_io_vec2_1),
    .io_vec2_2(VectorMul_7_io_vec2_2),
    .io_vec2_3(VectorMul_7_io_vec2_3),
    .io_vec2_4(VectorMul_7_io_vec2_4),
    .io_vec2_5(VectorMul_7_io_vec2_5),
    .io_vec2_6(VectorMul_7_io_vec2_6),
    .io_vec2_7(VectorMul_7_io_vec2_7),
    .io_vec2_8(VectorMul_7_io_vec2_8),
    .io_out(VectorMul_7_io_out)
  );
  VectorMul VectorMul_8 (
    .clock(VectorMul_8_clock),
    .reset(VectorMul_8_reset),
    .io_vec1_0(VectorMul_8_io_vec1_0),
    .io_vec1_1(VectorMul_8_io_vec1_1),
    .io_vec1_2(VectorMul_8_io_vec1_2),
    .io_vec1_3(VectorMul_8_io_vec1_3),
    .io_vec1_4(VectorMul_8_io_vec1_4),
    .io_vec1_5(VectorMul_8_io_vec1_5),
    .io_vec1_6(VectorMul_8_io_vec1_6),
    .io_vec1_7(VectorMul_8_io_vec1_7),
    .io_vec1_8(VectorMul_8_io_vec1_8),
    .io_vec2_0(VectorMul_8_io_vec2_0),
    .io_vec2_1(VectorMul_8_io_vec2_1),
    .io_vec2_2(VectorMul_8_io_vec2_2),
    .io_vec2_3(VectorMul_8_io_vec2_3),
    .io_vec2_4(VectorMul_8_io_vec2_4),
    .io_vec2_5(VectorMul_8_io_vec2_5),
    .io_vec2_6(VectorMul_8_io_vec2_6),
    .io_vec2_7(VectorMul_8_io_vec2_7),
    .io_vec2_8(VectorMul_8_io_vec2_8),
    .io_out(VectorMul_8_io_out)
  );
  VectorMul VectorMul_9 (
    .clock(VectorMul_9_clock),
    .reset(VectorMul_9_reset),
    .io_vec1_0(VectorMul_9_io_vec1_0),
    .io_vec1_1(VectorMul_9_io_vec1_1),
    .io_vec1_2(VectorMul_9_io_vec1_2),
    .io_vec1_3(VectorMul_9_io_vec1_3),
    .io_vec1_4(VectorMul_9_io_vec1_4),
    .io_vec1_5(VectorMul_9_io_vec1_5),
    .io_vec1_6(VectorMul_9_io_vec1_6),
    .io_vec1_7(VectorMul_9_io_vec1_7),
    .io_vec1_8(VectorMul_9_io_vec1_8),
    .io_vec2_0(VectorMul_9_io_vec2_0),
    .io_vec2_1(VectorMul_9_io_vec2_1),
    .io_vec2_2(VectorMul_9_io_vec2_2),
    .io_vec2_3(VectorMul_9_io_vec2_3),
    .io_vec2_4(VectorMul_9_io_vec2_4),
    .io_vec2_5(VectorMul_9_io_vec2_5),
    .io_vec2_6(VectorMul_9_io_vec2_6),
    .io_vec2_7(VectorMul_9_io_vec2_7),
    .io_vec2_8(VectorMul_9_io_vec2_8),
    .io_out(VectorMul_9_io_out)
  );
  VectorMul VectorMul_10 (
    .clock(VectorMul_10_clock),
    .reset(VectorMul_10_reset),
    .io_vec1_0(VectorMul_10_io_vec1_0),
    .io_vec1_1(VectorMul_10_io_vec1_1),
    .io_vec1_2(VectorMul_10_io_vec1_2),
    .io_vec1_3(VectorMul_10_io_vec1_3),
    .io_vec1_4(VectorMul_10_io_vec1_4),
    .io_vec1_5(VectorMul_10_io_vec1_5),
    .io_vec1_6(VectorMul_10_io_vec1_6),
    .io_vec1_7(VectorMul_10_io_vec1_7),
    .io_vec1_8(VectorMul_10_io_vec1_8),
    .io_vec2_0(VectorMul_10_io_vec2_0),
    .io_vec2_1(VectorMul_10_io_vec2_1),
    .io_vec2_2(VectorMul_10_io_vec2_2),
    .io_vec2_3(VectorMul_10_io_vec2_3),
    .io_vec2_4(VectorMul_10_io_vec2_4),
    .io_vec2_5(VectorMul_10_io_vec2_5),
    .io_vec2_6(VectorMul_10_io_vec2_6),
    .io_vec2_7(VectorMul_10_io_vec2_7),
    .io_vec2_8(VectorMul_10_io_vec2_8),
    .io_out(VectorMul_10_io_out)
  );
  VectorMul VectorMul_11 (
    .clock(VectorMul_11_clock),
    .reset(VectorMul_11_reset),
    .io_vec1_0(VectorMul_11_io_vec1_0),
    .io_vec1_1(VectorMul_11_io_vec1_1),
    .io_vec1_2(VectorMul_11_io_vec1_2),
    .io_vec1_3(VectorMul_11_io_vec1_3),
    .io_vec1_4(VectorMul_11_io_vec1_4),
    .io_vec1_5(VectorMul_11_io_vec1_5),
    .io_vec1_6(VectorMul_11_io_vec1_6),
    .io_vec1_7(VectorMul_11_io_vec1_7),
    .io_vec1_8(VectorMul_11_io_vec1_8),
    .io_vec2_0(VectorMul_11_io_vec2_0),
    .io_vec2_1(VectorMul_11_io_vec2_1),
    .io_vec2_2(VectorMul_11_io_vec2_2),
    .io_vec2_3(VectorMul_11_io_vec2_3),
    .io_vec2_4(VectorMul_11_io_vec2_4),
    .io_vec2_5(VectorMul_11_io_vec2_5),
    .io_vec2_6(VectorMul_11_io_vec2_6),
    .io_vec2_7(VectorMul_11_io_vec2_7),
    .io_vec2_8(VectorMul_11_io_vec2_8),
    .io_out(VectorMul_11_io_out)
  );
  VectorMul VectorMul_12 (
    .clock(VectorMul_12_clock),
    .reset(VectorMul_12_reset),
    .io_vec1_0(VectorMul_12_io_vec1_0),
    .io_vec1_1(VectorMul_12_io_vec1_1),
    .io_vec1_2(VectorMul_12_io_vec1_2),
    .io_vec1_3(VectorMul_12_io_vec1_3),
    .io_vec1_4(VectorMul_12_io_vec1_4),
    .io_vec1_5(VectorMul_12_io_vec1_5),
    .io_vec1_6(VectorMul_12_io_vec1_6),
    .io_vec1_7(VectorMul_12_io_vec1_7),
    .io_vec1_8(VectorMul_12_io_vec1_8),
    .io_vec2_0(VectorMul_12_io_vec2_0),
    .io_vec2_1(VectorMul_12_io_vec2_1),
    .io_vec2_2(VectorMul_12_io_vec2_2),
    .io_vec2_3(VectorMul_12_io_vec2_3),
    .io_vec2_4(VectorMul_12_io_vec2_4),
    .io_vec2_5(VectorMul_12_io_vec2_5),
    .io_vec2_6(VectorMul_12_io_vec2_6),
    .io_vec2_7(VectorMul_12_io_vec2_7),
    .io_vec2_8(VectorMul_12_io_vec2_8),
    .io_out(VectorMul_12_io_out)
  );
  VectorMul VectorMul_13 (
    .clock(VectorMul_13_clock),
    .reset(VectorMul_13_reset),
    .io_vec1_0(VectorMul_13_io_vec1_0),
    .io_vec1_1(VectorMul_13_io_vec1_1),
    .io_vec1_2(VectorMul_13_io_vec1_2),
    .io_vec1_3(VectorMul_13_io_vec1_3),
    .io_vec1_4(VectorMul_13_io_vec1_4),
    .io_vec1_5(VectorMul_13_io_vec1_5),
    .io_vec1_6(VectorMul_13_io_vec1_6),
    .io_vec1_7(VectorMul_13_io_vec1_7),
    .io_vec1_8(VectorMul_13_io_vec1_8),
    .io_vec2_0(VectorMul_13_io_vec2_0),
    .io_vec2_1(VectorMul_13_io_vec2_1),
    .io_vec2_2(VectorMul_13_io_vec2_2),
    .io_vec2_3(VectorMul_13_io_vec2_3),
    .io_vec2_4(VectorMul_13_io_vec2_4),
    .io_vec2_5(VectorMul_13_io_vec2_5),
    .io_vec2_6(VectorMul_13_io_vec2_6),
    .io_vec2_7(VectorMul_13_io_vec2_7),
    .io_vec2_8(VectorMul_13_io_vec2_8),
    .io_out(VectorMul_13_io_out)
  );
  VectorMul VectorMul_14 (
    .clock(VectorMul_14_clock),
    .reset(VectorMul_14_reset),
    .io_vec1_0(VectorMul_14_io_vec1_0),
    .io_vec1_1(VectorMul_14_io_vec1_1),
    .io_vec1_2(VectorMul_14_io_vec1_2),
    .io_vec1_3(VectorMul_14_io_vec1_3),
    .io_vec1_4(VectorMul_14_io_vec1_4),
    .io_vec1_5(VectorMul_14_io_vec1_5),
    .io_vec1_6(VectorMul_14_io_vec1_6),
    .io_vec1_7(VectorMul_14_io_vec1_7),
    .io_vec1_8(VectorMul_14_io_vec1_8),
    .io_vec2_0(VectorMul_14_io_vec2_0),
    .io_vec2_1(VectorMul_14_io_vec2_1),
    .io_vec2_2(VectorMul_14_io_vec2_2),
    .io_vec2_3(VectorMul_14_io_vec2_3),
    .io_vec2_4(VectorMul_14_io_vec2_4),
    .io_vec2_5(VectorMul_14_io_vec2_5),
    .io_vec2_6(VectorMul_14_io_vec2_6),
    .io_vec2_7(VectorMul_14_io_vec2_7),
    .io_vec2_8(VectorMul_14_io_vec2_8),
    .io_out(VectorMul_14_io_out)
  );
  VectorMul VectorMul_15 (
    .clock(VectorMul_15_clock),
    .reset(VectorMul_15_reset),
    .io_vec1_0(VectorMul_15_io_vec1_0),
    .io_vec1_1(VectorMul_15_io_vec1_1),
    .io_vec1_2(VectorMul_15_io_vec1_2),
    .io_vec1_3(VectorMul_15_io_vec1_3),
    .io_vec1_4(VectorMul_15_io_vec1_4),
    .io_vec1_5(VectorMul_15_io_vec1_5),
    .io_vec1_6(VectorMul_15_io_vec1_6),
    .io_vec1_7(VectorMul_15_io_vec1_7),
    .io_vec1_8(VectorMul_15_io_vec1_8),
    .io_vec2_0(VectorMul_15_io_vec2_0),
    .io_vec2_1(VectorMul_15_io_vec2_1),
    .io_vec2_2(VectorMul_15_io_vec2_2),
    .io_vec2_3(VectorMul_15_io_vec2_3),
    .io_vec2_4(VectorMul_15_io_vec2_4),
    .io_vec2_5(VectorMul_15_io_vec2_5),
    .io_vec2_6(VectorMul_15_io_vec2_6),
    .io_vec2_7(VectorMul_15_io_vec2_7),
    .io_vec2_8(VectorMul_15_io_vec2_8),
    .io_out(VectorMul_15_io_out)
  );
  VectorMul VectorMul_16 (
    .clock(VectorMul_16_clock),
    .reset(VectorMul_16_reset),
    .io_vec1_0(VectorMul_16_io_vec1_0),
    .io_vec1_1(VectorMul_16_io_vec1_1),
    .io_vec1_2(VectorMul_16_io_vec1_2),
    .io_vec1_3(VectorMul_16_io_vec1_3),
    .io_vec1_4(VectorMul_16_io_vec1_4),
    .io_vec1_5(VectorMul_16_io_vec1_5),
    .io_vec1_6(VectorMul_16_io_vec1_6),
    .io_vec1_7(VectorMul_16_io_vec1_7),
    .io_vec1_8(VectorMul_16_io_vec1_8),
    .io_vec2_0(VectorMul_16_io_vec2_0),
    .io_vec2_1(VectorMul_16_io_vec2_1),
    .io_vec2_2(VectorMul_16_io_vec2_2),
    .io_vec2_3(VectorMul_16_io_vec2_3),
    .io_vec2_4(VectorMul_16_io_vec2_4),
    .io_vec2_5(VectorMul_16_io_vec2_5),
    .io_vec2_6(VectorMul_16_io_vec2_6),
    .io_vec2_7(VectorMul_16_io_vec2_7),
    .io_vec2_8(VectorMul_16_io_vec2_8),
    .io_out(VectorMul_16_io_out)
  );
  VectorMul VectorMul_17 (
    .clock(VectorMul_17_clock),
    .reset(VectorMul_17_reset),
    .io_vec1_0(VectorMul_17_io_vec1_0),
    .io_vec1_1(VectorMul_17_io_vec1_1),
    .io_vec1_2(VectorMul_17_io_vec1_2),
    .io_vec1_3(VectorMul_17_io_vec1_3),
    .io_vec1_4(VectorMul_17_io_vec1_4),
    .io_vec1_5(VectorMul_17_io_vec1_5),
    .io_vec1_6(VectorMul_17_io_vec1_6),
    .io_vec1_7(VectorMul_17_io_vec1_7),
    .io_vec1_8(VectorMul_17_io_vec1_8),
    .io_vec2_0(VectorMul_17_io_vec2_0),
    .io_vec2_1(VectorMul_17_io_vec2_1),
    .io_vec2_2(VectorMul_17_io_vec2_2),
    .io_vec2_3(VectorMul_17_io_vec2_3),
    .io_vec2_4(VectorMul_17_io_vec2_4),
    .io_vec2_5(VectorMul_17_io_vec2_5),
    .io_vec2_6(VectorMul_17_io_vec2_6),
    .io_vec2_7(VectorMul_17_io_vec2_7),
    .io_vec2_8(VectorMul_17_io_vec2_8),
    .io_out(VectorMul_17_io_out)
  );
  VectorMul VectorMul_18 (
    .clock(VectorMul_18_clock),
    .reset(VectorMul_18_reset),
    .io_vec1_0(VectorMul_18_io_vec1_0),
    .io_vec1_1(VectorMul_18_io_vec1_1),
    .io_vec1_2(VectorMul_18_io_vec1_2),
    .io_vec1_3(VectorMul_18_io_vec1_3),
    .io_vec1_4(VectorMul_18_io_vec1_4),
    .io_vec1_5(VectorMul_18_io_vec1_5),
    .io_vec1_6(VectorMul_18_io_vec1_6),
    .io_vec1_7(VectorMul_18_io_vec1_7),
    .io_vec1_8(VectorMul_18_io_vec1_8),
    .io_vec2_0(VectorMul_18_io_vec2_0),
    .io_vec2_1(VectorMul_18_io_vec2_1),
    .io_vec2_2(VectorMul_18_io_vec2_2),
    .io_vec2_3(VectorMul_18_io_vec2_3),
    .io_vec2_4(VectorMul_18_io_vec2_4),
    .io_vec2_5(VectorMul_18_io_vec2_5),
    .io_vec2_6(VectorMul_18_io_vec2_6),
    .io_vec2_7(VectorMul_18_io_vec2_7),
    .io_vec2_8(VectorMul_18_io_vec2_8),
    .io_out(VectorMul_18_io_out)
  );
  VectorMul VectorMul_19 (
    .clock(VectorMul_19_clock),
    .reset(VectorMul_19_reset),
    .io_vec1_0(VectorMul_19_io_vec1_0),
    .io_vec1_1(VectorMul_19_io_vec1_1),
    .io_vec1_2(VectorMul_19_io_vec1_2),
    .io_vec1_3(VectorMul_19_io_vec1_3),
    .io_vec1_4(VectorMul_19_io_vec1_4),
    .io_vec1_5(VectorMul_19_io_vec1_5),
    .io_vec1_6(VectorMul_19_io_vec1_6),
    .io_vec1_7(VectorMul_19_io_vec1_7),
    .io_vec1_8(VectorMul_19_io_vec1_8),
    .io_vec2_0(VectorMul_19_io_vec2_0),
    .io_vec2_1(VectorMul_19_io_vec2_1),
    .io_vec2_2(VectorMul_19_io_vec2_2),
    .io_vec2_3(VectorMul_19_io_vec2_3),
    .io_vec2_4(VectorMul_19_io_vec2_4),
    .io_vec2_5(VectorMul_19_io_vec2_5),
    .io_vec2_6(VectorMul_19_io_vec2_6),
    .io_vec2_7(VectorMul_19_io_vec2_7),
    .io_vec2_8(VectorMul_19_io_vec2_8),
    .io_out(VectorMul_19_io_out)
  );
  VectorMul VectorMul_20 (
    .clock(VectorMul_20_clock),
    .reset(VectorMul_20_reset),
    .io_vec1_0(VectorMul_20_io_vec1_0),
    .io_vec1_1(VectorMul_20_io_vec1_1),
    .io_vec1_2(VectorMul_20_io_vec1_2),
    .io_vec1_3(VectorMul_20_io_vec1_3),
    .io_vec1_4(VectorMul_20_io_vec1_4),
    .io_vec1_5(VectorMul_20_io_vec1_5),
    .io_vec1_6(VectorMul_20_io_vec1_6),
    .io_vec1_7(VectorMul_20_io_vec1_7),
    .io_vec1_8(VectorMul_20_io_vec1_8),
    .io_vec2_0(VectorMul_20_io_vec2_0),
    .io_vec2_1(VectorMul_20_io_vec2_1),
    .io_vec2_2(VectorMul_20_io_vec2_2),
    .io_vec2_3(VectorMul_20_io_vec2_3),
    .io_vec2_4(VectorMul_20_io_vec2_4),
    .io_vec2_5(VectorMul_20_io_vec2_5),
    .io_vec2_6(VectorMul_20_io_vec2_6),
    .io_vec2_7(VectorMul_20_io_vec2_7),
    .io_vec2_8(VectorMul_20_io_vec2_8),
    .io_out(VectorMul_20_io_out)
  );
  VectorMul VectorMul_21 (
    .clock(VectorMul_21_clock),
    .reset(VectorMul_21_reset),
    .io_vec1_0(VectorMul_21_io_vec1_0),
    .io_vec1_1(VectorMul_21_io_vec1_1),
    .io_vec1_2(VectorMul_21_io_vec1_2),
    .io_vec1_3(VectorMul_21_io_vec1_3),
    .io_vec1_4(VectorMul_21_io_vec1_4),
    .io_vec1_5(VectorMul_21_io_vec1_5),
    .io_vec1_6(VectorMul_21_io_vec1_6),
    .io_vec1_7(VectorMul_21_io_vec1_7),
    .io_vec1_8(VectorMul_21_io_vec1_8),
    .io_vec2_0(VectorMul_21_io_vec2_0),
    .io_vec2_1(VectorMul_21_io_vec2_1),
    .io_vec2_2(VectorMul_21_io_vec2_2),
    .io_vec2_3(VectorMul_21_io_vec2_3),
    .io_vec2_4(VectorMul_21_io_vec2_4),
    .io_vec2_5(VectorMul_21_io_vec2_5),
    .io_vec2_6(VectorMul_21_io_vec2_6),
    .io_vec2_7(VectorMul_21_io_vec2_7),
    .io_vec2_8(VectorMul_21_io_vec2_8),
    .io_out(VectorMul_21_io_out)
  );
  VectorMul VectorMul_22 (
    .clock(VectorMul_22_clock),
    .reset(VectorMul_22_reset),
    .io_vec1_0(VectorMul_22_io_vec1_0),
    .io_vec1_1(VectorMul_22_io_vec1_1),
    .io_vec1_2(VectorMul_22_io_vec1_2),
    .io_vec1_3(VectorMul_22_io_vec1_3),
    .io_vec1_4(VectorMul_22_io_vec1_4),
    .io_vec1_5(VectorMul_22_io_vec1_5),
    .io_vec1_6(VectorMul_22_io_vec1_6),
    .io_vec1_7(VectorMul_22_io_vec1_7),
    .io_vec1_8(VectorMul_22_io_vec1_8),
    .io_vec2_0(VectorMul_22_io_vec2_0),
    .io_vec2_1(VectorMul_22_io_vec2_1),
    .io_vec2_2(VectorMul_22_io_vec2_2),
    .io_vec2_3(VectorMul_22_io_vec2_3),
    .io_vec2_4(VectorMul_22_io_vec2_4),
    .io_vec2_5(VectorMul_22_io_vec2_5),
    .io_vec2_6(VectorMul_22_io_vec2_6),
    .io_vec2_7(VectorMul_22_io_vec2_7),
    .io_vec2_8(VectorMul_22_io_vec2_8),
    .io_out(VectorMul_22_io_out)
  );
  VectorMul VectorMul_23 (
    .clock(VectorMul_23_clock),
    .reset(VectorMul_23_reset),
    .io_vec1_0(VectorMul_23_io_vec1_0),
    .io_vec1_1(VectorMul_23_io_vec1_1),
    .io_vec1_2(VectorMul_23_io_vec1_2),
    .io_vec1_3(VectorMul_23_io_vec1_3),
    .io_vec1_4(VectorMul_23_io_vec1_4),
    .io_vec1_5(VectorMul_23_io_vec1_5),
    .io_vec1_6(VectorMul_23_io_vec1_6),
    .io_vec1_7(VectorMul_23_io_vec1_7),
    .io_vec1_8(VectorMul_23_io_vec1_8),
    .io_vec2_0(VectorMul_23_io_vec2_0),
    .io_vec2_1(VectorMul_23_io_vec2_1),
    .io_vec2_2(VectorMul_23_io_vec2_2),
    .io_vec2_3(VectorMul_23_io_vec2_3),
    .io_vec2_4(VectorMul_23_io_vec2_4),
    .io_vec2_5(VectorMul_23_io_vec2_5),
    .io_vec2_6(VectorMul_23_io_vec2_6),
    .io_vec2_7(VectorMul_23_io_vec2_7),
    .io_vec2_8(VectorMul_23_io_vec2_8),
    .io_out(VectorMul_23_io_out)
  );
  VectorMul VectorMul_24 (
    .clock(VectorMul_24_clock),
    .reset(VectorMul_24_reset),
    .io_vec1_0(VectorMul_24_io_vec1_0),
    .io_vec1_1(VectorMul_24_io_vec1_1),
    .io_vec1_2(VectorMul_24_io_vec1_2),
    .io_vec1_3(VectorMul_24_io_vec1_3),
    .io_vec1_4(VectorMul_24_io_vec1_4),
    .io_vec1_5(VectorMul_24_io_vec1_5),
    .io_vec1_6(VectorMul_24_io_vec1_6),
    .io_vec1_7(VectorMul_24_io_vec1_7),
    .io_vec1_8(VectorMul_24_io_vec1_8),
    .io_vec2_0(VectorMul_24_io_vec2_0),
    .io_vec2_1(VectorMul_24_io_vec2_1),
    .io_vec2_2(VectorMul_24_io_vec2_2),
    .io_vec2_3(VectorMul_24_io_vec2_3),
    .io_vec2_4(VectorMul_24_io_vec2_4),
    .io_vec2_5(VectorMul_24_io_vec2_5),
    .io_vec2_6(VectorMul_24_io_vec2_6),
    .io_vec2_7(VectorMul_24_io_vec2_7),
    .io_vec2_8(VectorMul_24_io_vec2_8),
    .io_out(VectorMul_24_io_out)
  );
  assign io_out_0 = {{2'd0}, result_0};
  assign io_out_1 = {{2'd0}, result_1};
  assign io_out_2 = {{2'd0}, result_2};
  assign io_out_3 = {{2'd0}, result_3};
  assign io_out_4 = {{2'd0}, result_4};
  assign io_out_5 = {{2'd0}, result_5};
  assign io_out_6 = {{2'd0}, result_6};
  assign io_out_7 = {{2'd0}, result_7};
  assign io_out_8 = {{2'd0}, result_8};
  assign io_out_9 = {{2'd0}, result_9};
  assign io_out_10 = {{2'd0}, result_10};
  assign io_out_11 = {{2'd0}, result_11};
  assign io_out_12 = {{2'd0}, result_12};
  assign io_out_13 = {{2'd0}, result_13};
  assign io_out_14 = {{2'd0}, result_14};
  assign io_out_15 = {{2'd0}, result_15};
  assign io_out_16 = {{2'd0}, result_16};
  assign io_out_17 = {{2'd0}, result_17};
  assign io_out_18 = {{2'd0}, result_18};
  assign io_out_19 = {{2'd0}, result_19};
  assign io_out_20 = {{2'd0}, result_20};
  assign io_out_21 = {{2'd0}, result_21};
  assign io_out_22 = {{2'd0}, result_22};
  assign io_out_23 = {{2'd0}, result_23};
  assign io_out_24 = {{2'd0}, result_24};
  assign VectorMul_io_vec1_0 = 2'h0;
  assign VectorMul_io_vec1_1 = 2'h0;
  assign VectorMul_io_vec1_2 = 2'h0;
  assign VectorMul_io_vec1_3 = 2'h0;
  assign VectorMul_io_vec1_4 = _T_507_4;
  assign VectorMul_io_vec1_5 = _T_507_5;
  assign VectorMul_io_vec1_6 = 2'h0;
  assign VectorMul_io_vec1_7 = _T_507_7;
  assign VectorMul_io_vec1_8 = _T_507_8;
  assign VectorMul_io_vec2_0 = io_weights_0;
  assign VectorMul_io_vec2_1 = io_weights_1;
  assign VectorMul_io_vec2_2 = io_weights_2;
  assign VectorMul_io_vec2_3 = io_weights_3;
  assign VectorMul_io_vec2_4 = io_weights_4;
  assign VectorMul_io_vec2_5 = io_weights_5;
  assign VectorMul_io_vec2_6 = io_weights_6;
  assign VectorMul_io_vec2_7 = io_weights_7;
  assign VectorMul_io_vec2_8 = io_weights_8;
  assign VectorMul_clock = clock;
  assign VectorMul_reset = reset;
  assign VectorMul_1_io_vec1_0 = 2'h0;
  assign VectorMul_1_io_vec1_1 = 2'h0;
  assign VectorMul_1_io_vec1_2 = 2'h0;
  assign VectorMul_1_io_vec1_3 = _T_892_3;
  assign VectorMul_1_io_vec1_4 = _T_892_4;
  assign VectorMul_1_io_vec1_5 = _T_892_5;
  assign VectorMul_1_io_vec1_6 = _T_892_6;
  assign VectorMul_1_io_vec1_7 = _T_892_7;
  assign VectorMul_1_io_vec1_8 = _T_892_8;
  assign VectorMul_1_io_vec2_0 = io_weights_0;
  assign VectorMul_1_io_vec2_1 = io_weights_1;
  assign VectorMul_1_io_vec2_2 = io_weights_2;
  assign VectorMul_1_io_vec2_3 = io_weights_3;
  assign VectorMul_1_io_vec2_4 = io_weights_4;
  assign VectorMul_1_io_vec2_5 = io_weights_5;
  assign VectorMul_1_io_vec2_6 = io_weights_6;
  assign VectorMul_1_io_vec2_7 = io_weights_7;
  assign VectorMul_1_io_vec2_8 = io_weights_8;
  assign VectorMul_1_clock = clock;
  assign VectorMul_1_reset = reset;
  assign VectorMul_2_io_vec1_0 = 2'h0;
  assign VectorMul_2_io_vec1_1 = 2'h0;
  assign VectorMul_2_io_vec1_2 = 2'h0;
  assign VectorMul_2_io_vec1_3 = _T_1277_3;
  assign VectorMul_2_io_vec1_4 = _T_1277_4;
  assign VectorMul_2_io_vec1_5 = _T_1277_5;
  assign VectorMul_2_io_vec1_6 = _T_1277_6;
  assign VectorMul_2_io_vec1_7 = _T_1277_7;
  assign VectorMul_2_io_vec1_8 = _T_1277_8;
  assign VectorMul_2_io_vec2_0 = io_weights_0;
  assign VectorMul_2_io_vec2_1 = io_weights_1;
  assign VectorMul_2_io_vec2_2 = io_weights_2;
  assign VectorMul_2_io_vec2_3 = io_weights_3;
  assign VectorMul_2_io_vec2_4 = io_weights_4;
  assign VectorMul_2_io_vec2_5 = io_weights_5;
  assign VectorMul_2_io_vec2_6 = io_weights_6;
  assign VectorMul_2_io_vec2_7 = io_weights_7;
  assign VectorMul_2_io_vec2_8 = io_weights_8;
  assign VectorMul_2_clock = clock;
  assign VectorMul_2_reset = reset;
  assign VectorMul_3_io_vec1_0 = 2'h0;
  assign VectorMul_3_io_vec1_1 = 2'h0;
  assign VectorMul_3_io_vec1_2 = 2'h0;
  assign VectorMul_3_io_vec1_3 = _T_1662_3;
  assign VectorMul_3_io_vec1_4 = _T_1662_4;
  assign VectorMul_3_io_vec1_5 = _T_1662_5;
  assign VectorMul_3_io_vec1_6 = _T_1662_6;
  assign VectorMul_3_io_vec1_7 = _T_1662_7;
  assign VectorMul_3_io_vec1_8 = _T_1662_8;
  assign VectorMul_3_io_vec2_0 = io_weights_0;
  assign VectorMul_3_io_vec2_1 = io_weights_1;
  assign VectorMul_3_io_vec2_2 = io_weights_2;
  assign VectorMul_3_io_vec2_3 = io_weights_3;
  assign VectorMul_3_io_vec2_4 = io_weights_4;
  assign VectorMul_3_io_vec2_5 = io_weights_5;
  assign VectorMul_3_io_vec2_6 = io_weights_6;
  assign VectorMul_3_io_vec2_7 = io_weights_7;
  assign VectorMul_3_io_vec2_8 = io_weights_8;
  assign VectorMul_3_clock = clock;
  assign VectorMul_3_reset = reset;
  assign VectorMul_4_io_vec1_0 = 2'h0;
  assign VectorMul_4_io_vec1_1 = 2'h0;
  assign VectorMul_4_io_vec1_2 = 2'h0;
  assign VectorMul_4_io_vec1_3 = _T_2047_3;
  assign VectorMul_4_io_vec1_4 = _T_2047_4;
  assign VectorMul_4_io_vec1_5 = 2'h0;
  assign VectorMul_4_io_vec1_6 = _T_2047_6;
  assign VectorMul_4_io_vec1_7 = _T_2047_7;
  assign VectorMul_4_io_vec1_8 = 2'h0;
  assign VectorMul_4_io_vec2_0 = io_weights_0;
  assign VectorMul_4_io_vec2_1 = io_weights_1;
  assign VectorMul_4_io_vec2_2 = io_weights_2;
  assign VectorMul_4_io_vec2_3 = io_weights_3;
  assign VectorMul_4_io_vec2_4 = io_weights_4;
  assign VectorMul_4_io_vec2_5 = io_weights_5;
  assign VectorMul_4_io_vec2_6 = io_weights_6;
  assign VectorMul_4_io_vec2_7 = io_weights_7;
  assign VectorMul_4_io_vec2_8 = io_weights_8;
  assign VectorMul_4_clock = clock;
  assign VectorMul_4_reset = reset;
  assign VectorMul_5_io_vec1_0 = 2'h0;
  assign VectorMul_5_io_vec1_1 = _T_584_1;
  assign VectorMul_5_io_vec1_2 = _T_584_2;
  assign VectorMul_5_io_vec1_3 = 2'h0;
  assign VectorMul_5_io_vec1_4 = _T_584_4;
  assign VectorMul_5_io_vec1_5 = _T_584_5;
  assign VectorMul_5_io_vec1_6 = 2'h0;
  assign VectorMul_5_io_vec1_7 = _T_584_7;
  assign VectorMul_5_io_vec1_8 = _T_584_8;
  assign VectorMul_5_io_vec2_0 = io_weights_0;
  assign VectorMul_5_io_vec2_1 = io_weights_1;
  assign VectorMul_5_io_vec2_2 = io_weights_2;
  assign VectorMul_5_io_vec2_3 = io_weights_3;
  assign VectorMul_5_io_vec2_4 = io_weights_4;
  assign VectorMul_5_io_vec2_5 = io_weights_5;
  assign VectorMul_5_io_vec2_6 = io_weights_6;
  assign VectorMul_5_io_vec2_7 = io_weights_7;
  assign VectorMul_5_io_vec2_8 = io_weights_8;
  assign VectorMul_5_clock = clock;
  assign VectorMul_5_reset = reset;
  assign VectorMul_6_io_vec1_0 = _T_969_0;
  assign VectorMul_6_io_vec1_1 = _T_969_1;
  assign VectorMul_6_io_vec1_2 = _T_969_2;
  assign VectorMul_6_io_vec1_3 = _T_969_3;
  assign VectorMul_6_io_vec1_4 = _T_969_4;
  assign VectorMul_6_io_vec1_5 = _T_969_5;
  assign VectorMul_6_io_vec1_6 = _T_969_6;
  assign VectorMul_6_io_vec1_7 = _T_969_7;
  assign VectorMul_6_io_vec1_8 = _T_969_8;
  assign VectorMul_6_io_vec2_0 = io_weights_0;
  assign VectorMul_6_io_vec2_1 = io_weights_1;
  assign VectorMul_6_io_vec2_2 = io_weights_2;
  assign VectorMul_6_io_vec2_3 = io_weights_3;
  assign VectorMul_6_io_vec2_4 = io_weights_4;
  assign VectorMul_6_io_vec2_5 = io_weights_5;
  assign VectorMul_6_io_vec2_6 = io_weights_6;
  assign VectorMul_6_io_vec2_7 = io_weights_7;
  assign VectorMul_6_io_vec2_8 = io_weights_8;
  assign VectorMul_6_clock = clock;
  assign VectorMul_6_reset = reset;
  assign VectorMul_7_io_vec1_0 = _T_1354_0;
  assign VectorMul_7_io_vec1_1 = _T_1354_1;
  assign VectorMul_7_io_vec1_2 = _T_1354_2;
  assign VectorMul_7_io_vec1_3 = _T_1354_3;
  assign VectorMul_7_io_vec1_4 = _T_1354_4;
  assign VectorMul_7_io_vec1_5 = _T_1354_5;
  assign VectorMul_7_io_vec1_6 = _T_1354_6;
  assign VectorMul_7_io_vec1_7 = _T_1354_7;
  assign VectorMul_7_io_vec1_8 = _T_1354_8;
  assign VectorMul_7_io_vec2_0 = io_weights_0;
  assign VectorMul_7_io_vec2_1 = io_weights_1;
  assign VectorMul_7_io_vec2_2 = io_weights_2;
  assign VectorMul_7_io_vec2_3 = io_weights_3;
  assign VectorMul_7_io_vec2_4 = io_weights_4;
  assign VectorMul_7_io_vec2_5 = io_weights_5;
  assign VectorMul_7_io_vec2_6 = io_weights_6;
  assign VectorMul_7_io_vec2_7 = io_weights_7;
  assign VectorMul_7_io_vec2_8 = io_weights_8;
  assign VectorMul_7_clock = clock;
  assign VectorMul_7_reset = reset;
  assign VectorMul_8_io_vec1_0 = _T_1739_0;
  assign VectorMul_8_io_vec1_1 = _T_1739_1;
  assign VectorMul_8_io_vec1_2 = _T_1739_2;
  assign VectorMul_8_io_vec1_3 = _T_1739_3;
  assign VectorMul_8_io_vec1_4 = _T_1739_4;
  assign VectorMul_8_io_vec1_5 = _T_1739_5;
  assign VectorMul_8_io_vec1_6 = _T_1739_6;
  assign VectorMul_8_io_vec1_7 = _T_1739_7;
  assign VectorMul_8_io_vec1_8 = _T_1739_8;
  assign VectorMul_8_io_vec2_0 = io_weights_0;
  assign VectorMul_8_io_vec2_1 = io_weights_1;
  assign VectorMul_8_io_vec2_2 = io_weights_2;
  assign VectorMul_8_io_vec2_3 = io_weights_3;
  assign VectorMul_8_io_vec2_4 = io_weights_4;
  assign VectorMul_8_io_vec2_5 = io_weights_5;
  assign VectorMul_8_io_vec2_6 = io_weights_6;
  assign VectorMul_8_io_vec2_7 = io_weights_7;
  assign VectorMul_8_io_vec2_8 = io_weights_8;
  assign VectorMul_8_clock = clock;
  assign VectorMul_8_reset = reset;
  assign VectorMul_9_io_vec1_0 = _T_2124_0;
  assign VectorMul_9_io_vec1_1 = _T_2124_1;
  assign VectorMul_9_io_vec1_2 = 2'h0;
  assign VectorMul_9_io_vec1_3 = _T_2124_3;
  assign VectorMul_9_io_vec1_4 = _T_2124_4;
  assign VectorMul_9_io_vec1_5 = 2'h0;
  assign VectorMul_9_io_vec1_6 = _T_2124_6;
  assign VectorMul_9_io_vec1_7 = _T_2124_7;
  assign VectorMul_9_io_vec1_8 = 2'h0;
  assign VectorMul_9_io_vec2_0 = io_weights_0;
  assign VectorMul_9_io_vec2_1 = io_weights_1;
  assign VectorMul_9_io_vec2_2 = io_weights_2;
  assign VectorMul_9_io_vec2_3 = io_weights_3;
  assign VectorMul_9_io_vec2_4 = io_weights_4;
  assign VectorMul_9_io_vec2_5 = io_weights_5;
  assign VectorMul_9_io_vec2_6 = io_weights_6;
  assign VectorMul_9_io_vec2_7 = io_weights_7;
  assign VectorMul_9_io_vec2_8 = io_weights_8;
  assign VectorMul_9_clock = clock;
  assign VectorMul_9_reset = reset;
  assign VectorMul_10_io_vec1_0 = 2'h0;
  assign VectorMul_10_io_vec1_1 = _T_661_1;
  assign VectorMul_10_io_vec1_2 = _T_661_2;
  assign VectorMul_10_io_vec1_3 = 2'h0;
  assign VectorMul_10_io_vec1_4 = _T_661_4;
  assign VectorMul_10_io_vec1_5 = _T_661_5;
  assign VectorMul_10_io_vec1_6 = 2'h0;
  assign VectorMul_10_io_vec1_7 = _T_661_7;
  assign VectorMul_10_io_vec1_8 = _T_661_8;
  assign VectorMul_10_io_vec2_0 = io_weights_0;
  assign VectorMul_10_io_vec2_1 = io_weights_1;
  assign VectorMul_10_io_vec2_2 = io_weights_2;
  assign VectorMul_10_io_vec2_3 = io_weights_3;
  assign VectorMul_10_io_vec2_4 = io_weights_4;
  assign VectorMul_10_io_vec2_5 = io_weights_5;
  assign VectorMul_10_io_vec2_6 = io_weights_6;
  assign VectorMul_10_io_vec2_7 = io_weights_7;
  assign VectorMul_10_io_vec2_8 = io_weights_8;
  assign VectorMul_10_clock = clock;
  assign VectorMul_10_reset = reset;
  assign VectorMul_11_io_vec1_0 = _T_1046_0;
  assign VectorMul_11_io_vec1_1 = _T_1046_1;
  assign VectorMul_11_io_vec1_2 = _T_1046_2;
  assign VectorMul_11_io_vec1_3 = _T_1046_3;
  assign VectorMul_11_io_vec1_4 = _T_1046_4;
  assign VectorMul_11_io_vec1_5 = _T_1046_5;
  assign VectorMul_11_io_vec1_6 = _T_1046_6;
  assign VectorMul_11_io_vec1_7 = _T_1046_7;
  assign VectorMul_11_io_vec1_8 = _T_1046_8;
  assign VectorMul_11_io_vec2_0 = io_weights_0;
  assign VectorMul_11_io_vec2_1 = io_weights_1;
  assign VectorMul_11_io_vec2_2 = io_weights_2;
  assign VectorMul_11_io_vec2_3 = io_weights_3;
  assign VectorMul_11_io_vec2_4 = io_weights_4;
  assign VectorMul_11_io_vec2_5 = io_weights_5;
  assign VectorMul_11_io_vec2_6 = io_weights_6;
  assign VectorMul_11_io_vec2_7 = io_weights_7;
  assign VectorMul_11_io_vec2_8 = io_weights_8;
  assign VectorMul_11_clock = clock;
  assign VectorMul_11_reset = reset;
  assign VectorMul_12_io_vec1_0 = _T_1431_0;
  assign VectorMul_12_io_vec1_1 = _T_1431_1;
  assign VectorMul_12_io_vec1_2 = _T_1431_2;
  assign VectorMul_12_io_vec1_3 = _T_1431_3;
  assign VectorMul_12_io_vec1_4 = _T_1431_4;
  assign VectorMul_12_io_vec1_5 = _T_1431_5;
  assign VectorMul_12_io_vec1_6 = _T_1431_6;
  assign VectorMul_12_io_vec1_7 = _T_1431_7;
  assign VectorMul_12_io_vec1_8 = _T_1431_8;
  assign VectorMul_12_io_vec2_0 = io_weights_0;
  assign VectorMul_12_io_vec2_1 = io_weights_1;
  assign VectorMul_12_io_vec2_2 = io_weights_2;
  assign VectorMul_12_io_vec2_3 = io_weights_3;
  assign VectorMul_12_io_vec2_4 = io_weights_4;
  assign VectorMul_12_io_vec2_5 = io_weights_5;
  assign VectorMul_12_io_vec2_6 = io_weights_6;
  assign VectorMul_12_io_vec2_7 = io_weights_7;
  assign VectorMul_12_io_vec2_8 = io_weights_8;
  assign VectorMul_12_clock = clock;
  assign VectorMul_12_reset = reset;
  assign VectorMul_13_io_vec1_0 = _T_1816_0;
  assign VectorMul_13_io_vec1_1 = _T_1816_1;
  assign VectorMul_13_io_vec1_2 = _T_1816_2;
  assign VectorMul_13_io_vec1_3 = _T_1816_3;
  assign VectorMul_13_io_vec1_4 = _T_1816_4;
  assign VectorMul_13_io_vec1_5 = _T_1816_5;
  assign VectorMul_13_io_vec1_6 = _T_1816_6;
  assign VectorMul_13_io_vec1_7 = _T_1816_7;
  assign VectorMul_13_io_vec1_8 = _T_1816_8;
  assign VectorMul_13_io_vec2_0 = io_weights_0;
  assign VectorMul_13_io_vec2_1 = io_weights_1;
  assign VectorMul_13_io_vec2_2 = io_weights_2;
  assign VectorMul_13_io_vec2_3 = io_weights_3;
  assign VectorMul_13_io_vec2_4 = io_weights_4;
  assign VectorMul_13_io_vec2_5 = io_weights_5;
  assign VectorMul_13_io_vec2_6 = io_weights_6;
  assign VectorMul_13_io_vec2_7 = io_weights_7;
  assign VectorMul_13_io_vec2_8 = io_weights_8;
  assign VectorMul_13_clock = clock;
  assign VectorMul_13_reset = reset;
  assign VectorMul_14_io_vec1_0 = _T_2201_0;
  assign VectorMul_14_io_vec1_1 = _T_2201_1;
  assign VectorMul_14_io_vec1_2 = 2'h0;
  assign VectorMul_14_io_vec1_3 = _T_2201_3;
  assign VectorMul_14_io_vec1_4 = _T_2201_4;
  assign VectorMul_14_io_vec1_5 = 2'h0;
  assign VectorMul_14_io_vec1_6 = _T_2201_6;
  assign VectorMul_14_io_vec1_7 = _T_2201_7;
  assign VectorMul_14_io_vec1_8 = 2'h0;
  assign VectorMul_14_io_vec2_0 = io_weights_0;
  assign VectorMul_14_io_vec2_1 = io_weights_1;
  assign VectorMul_14_io_vec2_2 = io_weights_2;
  assign VectorMul_14_io_vec2_3 = io_weights_3;
  assign VectorMul_14_io_vec2_4 = io_weights_4;
  assign VectorMul_14_io_vec2_5 = io_weights_5;
  assign VectorMul_14_io_vec2_6 = io_weights_6;
  assign VectorMul_14_io_vec2_7 = io_weights_7;
  assign VectorMul_14_io_vec2_8 = io_weights_8;
  assign VectorMul_14_clock = clock;
  assign VectorMul_14_reset = reset;
  assign VectorMul_15_io_vec1_0 = 2'h0;
  assign VectorMul_15_io_vec1_1 = _T_738_1;
  assign VectorMul_15_io_vec1_2 = _T_738_2;
  assign VectorMul_15_io_vec1_3 = 2'h0;
  assign VectorMul_15_io_vec1_4 = _T_738_4;
  assign VectorMul_15_io_vec1_5 = _T_738_5;
  assign VectorMul_15_io_vec1_6 = 2'h0;
  assign VectorMul_15_io_vec1_7 = _T_738_7;
  assign VectorMul_15_io_vec1_8 = _T_738_8;
  assign VectorMul_15_io_vec2_0 = io_weights_0;
  assign VectorMul_15_io_vec2_1 = io_weights_1;
  assign VectorMul_15_io_vec2_2 = io_weights_2;
  assign VectorMul_15_io_vec2_3 = io_weights_3;
  assign VectorMul_15_io_vec2_4 = io_weights_4;
  assign VectorMul_15_io_vec2_5 = io_weights_5;
  assign VectorMul_15_io_vec2_6 = io_weights_6;
  assign VectorMul_15_io_vec2_7 = io_weights_7;
  assign VectorMul_15_io_vec2_8 = io_weights_8;
  assign VectorMul_15_clock = clock;
  assign VectorMul_15_reset = reset;
  assign VectorMul_16_io_vec1_0 = _T_1123_0;
  assign VectorMul_16_io_vec1_1 = _T_1123_1;
  assign VectorMul_16_io_vec1_2 = _T_1123_2;
  assign VectorMul_16_io_vec1_3 = _T_1123_3;
  assign VectorMul_16_io_vec1_4 = _T_1123_4;
  assign VectorMul_16_io_vec1_5 = _T_1123_5;
  assign VectorMul_16_io_vec1_6 = _T_1123_6;
  assign VectorMul_16_io_vec1_7 = _T_1123_7;
  assign VectorMul_16_io_vec1_8 = _T_1123_8;
  assign VectorMul_16_io_vec2_0 = io_weights_0;
  assign VectorMul_16_io_vec2_1 = io_weights_1;
  assign VectorMul_16_io_vec2_2 = io_weights_2;
  assign VectorMul_16_io_vec2_3 = io_weights_3;
  assign VectorMul_16_io_vec2_4 = io_weights_4;
  assign VectorMul_16_io_vec2_5 = io_weights_5;
  assign VectorMul_16_io_vec2_6 = io_weights_6;
  assign VectorMul_16_io_vec2_7 = io_weights_7;
  assign VectorMul_16_io_vec2_8 = io_weights_8;
  assign VectorMul_16_clock = clock;
  assign VectorMul_16_reset = reset;
  assign VectorMul_17_io_vec1_0 = _T_1508_0;
  assign VectorMul_17_io_vec1_1 = _T_1508_1;
  assign VectorMul_17_io_vec1_2 = _T_1508_2;
  assign VectorMul_17_io_vec1_3 = _T_1508_3;
  assign VectorMul_17_io_vec1_4 = _T_1508_4;
  assign VectorMul_17_io_vec1_5 = _T_1508_5;
  assign VectorMul_17_io_vec1_6 = _T_1508_6;
  assign VectorMul_17_io_vec1_7 = _T_1508_7;
  assign VectorMul_17_io_vec1_8 = _T_1508_8;
  assign VectorMul_17_io_vec2_0 = io_weights_0;
  assign VectorMul_17_io_vec2_1 = io_weights_1;
  assign VectorMul_17_io_vec2_2 = io_weights_2;
  assign VectorMul_17_io_vec2_3 = io_weights_3;
  assign VectorMul_17_io_vec2_4 = io_weights_4;
  assign VectorMul_17_io_vec2_5 = io_weights_5;
  assign VectorMul_17_io_vec2_6 = io_weights_6;
  assign VectorMul_17_io_vec2_7 = io_weights_7;
  assign VectorMul_17_io_vec2_8 = io_weights_8;
  assign VectorMul_17_clock = clock;
  assign VectorMul_17_reset = reset;
  assign VectorMul_18_io_vec1_0 = _T_1893_0;
  assign VectorMul_18_io_vec1_1 = _T_1893_1;
  assign VectorMul_18_io_vec1_2 = _T_1893_2;
  assign VectorMul_18_io_vec1_3 = _T_1893_3;
  assign VectorMul_18_io_vec1_4 = _T_1893_4;
  assign VectorMul_18_io_vec1_5 = _T_1893_5;
  assign VectorMul_18_io_vec1_6 = _T_1893_6;
  assign VectorMul_18_io_vec1_7 = _T_1893_7;
  assign VectorMul_18_io_vec1_8 = _T_1893_8;
  assign VectorMul_18_io_vec2_0 = io_weights_0;
  assign VectorMul_18_io_vec2_1 = io_weights_1;
  assign VectorMul_18_io_vec2_2 = io_weights_2;
  assign VectorMul_18_io_vec2_3 = io_weights_3;
  assign VectorMul_18_io_vec2_4 = io_weights_4;
  assign VectorMul_18_io_vec2_5 = io_weights_5;
  assign VectorMul_18_io_vec2_6 = io_weights_6;
  assign VectorMul_18_io_vec2_7 = io_weights_7;
  assign VectorMul_18_io_vec2_8 = io_weights_8;
  assign VectorMul_18_clock = clock;
  assign VectorMul_18_reset = reset;
  assign VectorMul_19_io_vec1_0 = _T_2278_0;
  assign VectorMul_19_io_vec1_1 = _T_2278_1;
  assign VectorMul_19_io_vec1_2 = 2'h0;
  assign VectorMul_19_io_vec1_3 = _T_2278_3;
  assign VectorMul_19_io_vec1_4 = _T_2278_4;
  assign VectorMul_19_io_vec1_5 = 2'h0;
  assign VectorMul_19_io_vec1_6 = _T_2278_6;
  assign VectorMul_19_io_vec1_7 = _T_2278_7;
  assign VectorMul_19_io_vec1_8 = 2'h0;
  assign VectorMul_19_io_vec2_0 = io_weights_0;
  assign VectorMul_19_io_vec2_1 = io_weights_1;
  assign VectorMul_19_io_vec2_2 = io_weights_2;
  assign VectorMul_19_io_vec2_3 = io_weights_3;
  assign VectorMul_19_io_vec2_4 = io_weights_4;
  assign VectorMul_19_io_vec2_5 = io_weights_5;
  assign VectorMul_19_io_vec2_6 = io_weights_6;
  assign VectorMul_19_io_vec2_7 = io_weights_7;
  assign VectorMul_19_io_vec2_8 = io_weights_8;
  assign VectorMul_19_clock = clock;
  assign VectorMul_19_reset = reset;
  assign VectorMul_20_io_vec1_0 = 2'h0;
  assign VectorMul_20_io_vec1_1 = _T_815_1;
  assign VectorMul_20_io_vec1_2 = _T_815_2;
  assign VectorMul_20_io_vec1_3 = 2'h0;
  assign VectorMul_20_io_vec1_4 = _T_815_4;
  assign VectorMul_20_io_vec1_5 = _T_815_5;
  assign VectorMul_20_io_vec1_6 = 2'h0;
  assign VectorMul_20_io_vec1_7 = 2'h0;
  assign VectorMul_20_io_vec1_8 = 2'h0;
  assign VectorMul_20_io_vec2_0 = io_weights_0;
  assign VectorMul_20_io_vec2_1 = io_weights_1;
  assign VectorMul_20_io_vec2_2 = io_weights_2;
  assign VectorMul_20_io_vec2_3 = io_weights_3;
  assign VectorMul_20_io_vec2_4 = io_weights_4;
  assign VectorMul_20_io_vec2_5 = io_weights_5;
  assign VectorMul_20_io_vec2_6 = io_weights_6;
  assign VectorMul_20_io_vec2_7 = io_weights_7;
  assign VectorMul_20_io_vec2_8 = io_weights_8;
  assign VectorMul_20_clock = clock;
  assign VectorMul_20_reset = reset;
  assign VectorMul_21_io_vec1_0 = _T_1200_0;
  assign VectorMul_21_io_vec1_1 = _T_1200_1;
  assign VectorMul_21_io_vec1_2 = _T_1200_2;
  assign VectorMul_21_io_vec1_3 = _T_1200_3;
  assign VectorMul_21_io_vec1_4 = _T_1200_4;
  assign VectorMul_21_io_vec1_5 = _T_1200_5;
  assign VectorMul_21_io_vec1_6 = 2'h0;
  assign VectorMul_21_io_vec1_7 = 2'h0;
  assign VectorMul_21_io_vec1_8 = 2'h0;
  assign VectorMul_21_io_vec2_0 = io_weights_0;
  assign VectorMul_21_io_vec2_1 = io_weights_1;
  assign VectorMul_21_io_vec2_2 = io_weights_2;
  assign VectorMul_21_io_vec2_3 = io_weights_3;
  assign VectorMul_21_io_vec2_4 = io_weights_4;
  assign VectorMul_21_io_vec2_5 = io_weights_5;
  assign VectorMul_21_io_vec2_6 = io_weights_6;
  assign VectorMul_21_io_vec2_7 = io_weights_7;
  assign VectorMul_21_io_vec2_8 = io_weights_8;
  assign VectorMul_21_clock = clock;
  assign VectorMul_21_reset = reset;
  assign VectorMul_22_io_vec1_0 = _T_1585_0;
  assign VectorMul_22_io_vec1_1 = _T_1585_1;
  assign VectorMul_22_io_vec1_2 = _T_1585_2;
  assign VectorMul_22_io_vec1_3 = _T_1585_3;
  assign VectorMul_22_io_vec1_4 = _T_1585_4;
  assign VectorMul_22_io_vec1_5 = _T_1585_5;
  assign VectorMul_22_io_vec1_6 = 2'h0;
  assign VectorMul_22_io_vec1_7 = 2'h0;
  assign VectorMul_22_io_vec1_8 = 2'h0;
  assign VectorMul_22_io_vec2_0 = io_weights_0;
  assign VectorMul_22_io_vec2_1 = io_weights_1;
  assign VectorMul_22_io_vec2_2 = io_weights_2;
  assign VectorMul_22_io_vec2_3 = io_weights_3;
  assign VectorMul_22_io_vec2_4 = io_weights_4;
  assign VectorMul_22_io_vec2_5 = io_weights_5;
  assign VectorMul_22_io_vec2_6 = io_weights_6;
  assign VectorMul_22_io_vec2_7 = io_weights_7;
  assign VectorMul_22_io_vec2_8 = io_weights_8;
  assign VectorMul_22_clock = clock;
  assign VectorMul_22_reset = reset;
  assign VectorMul_23_io_vec1_0 = _T_1970_0;
  assign VectorMul_23_io_vec1_1 = _T_1970_1;
  assign VectorMul_23_io_vec1_2 = _T_1970_2;
  assign VectorMul_23_io_vec1_3 = _T_1970_3;
  assign VectorMul_23_io_vec1_4 = _T_1970_4;
  assign VectorMul_23_io_vec1_5 = _T_1970_5;
  assign VectorMul_23_io_vec1_6 = 2'h0;
  assign VectorMul_23_io_vec1_7 = 2'h0;
  assign VectorMul_23_io_vec1_8 = 2'h0;
  assign VectorMul_23_io_vec2_0 = io_weights_0;
  assign VectorMul_23_io_vec2_1 = io_weights_1;
  assign VectorMul_23_io_vec2_2 = io_weights_2;
  assign VectorMul_23_io_vec2_3 = io_weights_3;
  assign VectorMul_23_io_vec2_4 = io_weights_4;
  assign VectorMul_23_io_vec2_5 = io_weights_5;
  assign VectorMul_23_io_vec2_6 = io_weights_6;
  assign VectorMul_23_io_vec2_7 = io_weights_7;
  assign VectorMul_23_io_vec2_8 = io_weights_8;
  assign VectorMul_23_clock = clock;
  assign VectorMul_23_reset = reset;
  assign VectorMul_24_io_vec1_0 = _T_2355_0;
  assign VectorMul_24_io_vec1_1 = _T_2355_1;
  assign VectorMul_24_io_vec1_2 = 2'h0;
  assign VectorMul_24_io_vec1_3 = _T_2355_3;
  assign VectorMul_24_io_vec1_4 = _T_2355_4;
  assign VectorMul_24_io_vec1_5 = 2'h0;
  assign VectorMul_24_io_vec1_6 = 2'h0;
  assign VectorMul_24_io_vec1_7 = 2'h0;
  assign VectorMul_24_io_vec1_8 = 2'h0;
  assign VectorMul_24_io_vec2_0 = io_weights_0;
  assign VectorMul_24_io_vec2_1 = io_weights_1;
  assign VectorMul_24_io_vec2_2 = io_weights_2;
  assign VectorMul_24_io_vec2_3 = io_weights_3;
  assign VectorMul_24_io_vec2_4 = io_weights_4;
  assign VectorMul_24_io_vec2_5 = io_weights_5;
  assign VectorMul_24_io_vec2_6 = io_weights_6;
  assign VectorMul_24_io_vec2_7 = io_weights_7;
  assign VectorMul_24_io_vec2_8 = io_weights_8;
  assign VectorMul_24_clock = clock;
  assign VectorMul_24_reset = reset;
  assign result_0 = VectorMul_io_out;
  assign result_1 = VectorMul_1_io_out;
  assign result_2 = VectorMul_2_io_out;
  assign result_3 = VectorMul_3_io_out;
  assign result_4 = VectorMul_4_io_out;
  assign result_5 = VectorMul_5_io_out;
  assign result_6 = VectorMul_6_io_out;
  assign result_7 = VectorMul_7_io_out;
  assign result_8 = VectorMul_8_io_out;
  assign result_9 = VectorMul_9_io_out;
  assign result_10 = VectorMul_10_io_out;
  assign result_11 = VectorMul_11_io_out;
  assign result_12 = VectorMul_12_io_out;
  assign result_13 = VectorMul_13_io_out;
  assign result_14 = VectorMul_14_io_out;
  assign result_15 = VectorMul_15_io_out;
  assign result_16 = VectorMul_16_io_out;
  assign result_17 = VectorMul_17_io_out;
  assign result_18 = VectorMul_18_io_out;
  assign result_19 = VectorMul_19_io_out;
  assign result_20 = VectorMul_20_io_out;
  assign result_21 = VectorMul_21_io_out;
  assign result_22 = VectorMul_22_io_out;
  assign result_23 = VectorMul_23_io_out;
  assign result_24 = VectorMul_24_io_out;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  xx_8 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  xx_9 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  xx_10 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  xx_11 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  xx_12 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  xx_15 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  xx_16 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  xx_17 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  xx_18 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  xx_19 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  xx_22 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  xx_23 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  xx_24 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  xx_25 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  xx_26 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  xx_29 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  xx_30 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  xx_31 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  xx_32 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  xx_33 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  xx_36 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  xx_37 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  xx_38 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  xx_39 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  xx_40 = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_507_4 = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_507_5 = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_507_7 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_507_8 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_584_1 = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_584_2 = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_584_4 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_584_5 = _RAND_32[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_584_7 = _RAND_33[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_584_8 = _RAND_34[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_661_1 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_661_2 = _RAND_36[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_661_4 = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_661_5 = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_661_7 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_661_8 = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_738_1 = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_738_2 = _RAND_42[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_738_4 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_738_5 = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_738_7 = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_738_8 = _RAND_46[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_815_1 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_815_2 = _RAND_48[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_815_4 = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_815_5 = _RAND_50[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_892_3 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_892_4 = _RAND_52[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_892_5 = _RAND_53[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_892_6 = _RAND_54[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_892_7 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_892_8 = _RAND_56[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_969_0 = _RAND_57[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_969_1 = _RAND_58[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_969_2 = _RAND_59[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_969_3 = _RAND_60[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_969_4 = _RAND_61[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_969_5 = _RAND_62[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_969_6 = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_969_7 = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_969_8 = _RAND_65[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_1046_0 = _RAND_66[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_1046_1 = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_1046_2 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_1046_3 = _RAND_69[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_1046_4 = _RAND_70[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_1046_5 = _RAND_71[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_1046_6 = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_1046_7 = _RAND_73[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_1046_8 = _RAND_74[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_1123_0 = _RAND_75[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_1123_1 = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_1123_2 = _RAND_77[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_1123_3 = _RAND_78[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_1123_4 = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_1123_5 = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_1123_6 = _RAND_81[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_1123_7 = _RAND_82[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_1123_8 = _RAND_83[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_1200_0 = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_1200_1 = _RAND_85[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_1200_2 = _RAND_86[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_1200_3 = _RAND_87[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_1200_4 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_1200_5 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_1277_3 = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_1277_4 = _RAND_91[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_1277_5 = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_1277_6 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_1277_7 = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_1277_8 = _RAND_95[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_1354_0 = _RAND_96[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_1354_1 = _RAND_97[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_1354_2 = _RAND_98[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_1354_3 = _RAND_99[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_1354_4 = _RAND_100[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_1354_5 = _RAND_101[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_1354_6 = _RAND_102[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_1354_7 = _RAND_103[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_1354_8 = _RAND_104[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_1431_0 = _RAND_105[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_1431_1 = _RAND_106[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_1431_2 = _RAND_107[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_1431_3 = _RAND_108[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_1431_4 = _RAND_109[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_1431_5 = _RAND_110[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_1431_6 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_1431_7 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_1431_8 = _RAND_113[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_1508_0 = _RAND_114[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_1508_1 = _RAND_115[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_1508_2 = _RAND_116[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_1508_3 = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_1508_4 = _RAND_118[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_1508_5 = _RAND_119[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_1508_6 = _RAND_120[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_1508_7 = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_1508_8 = _RAND_122[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_1585_0 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_1585_1 = _RAND_124[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_1585_2 = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_1585_3 = _RAND_126[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_1585_4 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_1585_5 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_1662_3 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_1662_4 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_1662_5 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_1662_6 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_1662_7 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_1662_8 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_1739_0 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_1739_1 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_1739_2 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_1739_3 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_1739_4 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_1739_5 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_1739_6 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_1739_7 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_1739_8 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_1816_0 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_1816_1 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_1816_2 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_1816_3 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_1816_4 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_1816_5 = _RAND_149[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_1816_6 = _RAND_150[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_1816_7 = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_1816_8 = _RAND_152[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_1893_0 = _RAND_153[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_1893_1 = _RAND_154[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_1893_2 = _RAND_155[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_1893_3 = _RAND_156[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_1893_4 = _RAND_157[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_1893_5 = _RAND_158[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_1893_6 = _RAND_159[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_1893_7 = _RAND_160[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_1893_8 = _RAND_161[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_1970_0 = _RAND_162[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_1970_1 = _RAND_163[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_1970_2 = _RAND_164[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_1970_3 = _RAND_165[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_1970_4 = _RAND_166[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_1970_5 = _RAND_167[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_2047_3 = _RAND_168[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_2047_4 = _RAND_169[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_2047_6 = _RAND_170[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_2047_7 = _RAND_171[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_2124_0 = _RAND_172[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_2124_1 = _RAND_173[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _T_2124_3 = _RAND_174[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _T_2124_4 = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _T_2124_6 = _RAND_176[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _T_2124_7 = _RAND_177[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _T_2201_0 = _RAND_178[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _T_2201_1 = _RAND_179[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  _T_2201_3 = _RAND_180[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  _T_2201_4 = _RAND_181[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  _T_2201_6 = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  _T_2201_7 = _RAND_183[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  _T_2278_0 = _RAND_184[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  _T_2278_1 = _RAND_185[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  _T_2278_3 = _RAND_186[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  _T_2278_4 = _RAND_187[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  _T_2278_6 = _RAND_188[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  _T_2278_7 = _RAND_189[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  _T_2355_0 = _RAND_190[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  _T_2355_1 = _RAND_191[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  _T_2355_3 = _RAND_192[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  _T_2355_4 = _RAND_193[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      xx_8 <= 2'h0;
    end else begin
      xx_8 <= io_mask_0;
    end
    if (reset) begin
      xx_9 <= 2'h0;
    end else begin
      xx_9 <= io_mask_1;
    end
    if (reset) begin
      xx_10 <= 2'h0;
    end else begin
      xx_10 <= io_mask_2;
    end
    if (reset) begin
      xx_11 <= 2'h0;
    end else begin
      xx_11 <= io_mask_3;
    end
    if (reset) begin
      xx_12 <= 2'h0;
    end else begin
      xx_12 <= io_mask_4;
    end
    if (reset) begin
      xx_15 <= 2'h0;
    end else begin
      xx_15 <= io_mask_5;
    end
    if (reset) begin
      xx_16 <= 2'h0;
    end else begin
      xx_16 <= io_mask_6;
    end
    if (reset) begin
      xx_17 <= 2'h0;
    end else begin
      xx_17 <= io_mask_7;
    end
    if (reset) begin
      xx_18 <= 2'h0;
    end else begin
      xx_18 <= io_mask_8;
    end
    if (reset) begin
      xx_19 <= 2'h0;
    end else begin
      xx_19 <= io_mask_9;
    end
    if (reset) begin
      xx_22 <= 2'h0;
    end else begin
      xx_22 <= io_mask_10;
    end
    if (reset) begin
      xx_23 <= 2'h0;
    end else begin
      xx_23 <= io_mask_11;
    end
    if (reset) begin
      xx_24 <= 2'h0;
    end else begin
      xx_24 <= io_mask_12;
    end
    if (reset) begin
      xx_25 <= 2'h0;
    end else begin
      xx_25 <= io_mask_13;
    end
    if (reset) begin
      xx_26 <= 2'h0;
    end else begin
      xx_26 <= io_mask_14;
    end
    if (reset) begin
      xx_29 <= 2'h0;
    end else begin
      xx_29 <= io_mask_15;
    end
    if (reset) begin
      xx_30 <= 2'h0;
    end else begin
      xx_30 <= io_mask_16;
    end
    if (reset) begin
      xx_31 <= 2'h0;
    end else begin
      xx_31 <= io_mask_17;
    end
    if (reset) begin
      xx_32 <= 2'h0;
    end else begin
      xx_32 <= io_mask_18;
    end
    if (reset) begin
      xx_33 <= 2'h0;
    end else begin
      xx_33 <= io_mask_19;
    end
    if (reset) begin
      xx_36 <= 2'h0;
    end else begin
      xx_36 <= io_mask_20;
    end
    if (reset) begin
      xx_37 <= 2'h0;
    end else begin
      xx_37 <= io_mask_21;
    end
    if (reset) begin
      xx_38 <= 2'h0;
    end else begin
      xx_38 <= io_mask_22;
    end
    if (reset) begin
      xx_39 <= 2'h0;
    end else begin
      xx_39 <= io_mask_23;
    end
    if (reset) begin
      xx_40 <= 2'h0;
    end else begin
      xx_40 <= io_mask_24;
    end
    if (reset) begin
      _T_507_4 <= 2'h0;
    end else begin
      _T_507_4 <= xx_8;
    end
    if (reset) begin
      _T_507_5 <= 2'h0;
    end else begin
      _T_507_5 <= xx_9;
    end
    if (reset) begin
      _T_507_7 <= 2'h0;
    end else begin
      _T_507_7 <= xx_15;
    end
    if (reset) begin
      _T_507_8 <= 2'h0;
    end else begin
      _T_507_8 <= xx_16;
    end
    if (reset) begin
      _T_584_1 <= 2'h0;
    end else begin
      _T_584_1 <= xx_8;
    end
    if (reset) begin
      _T_584_2 <= 2'h0;
    end else begin
      _T_584_2 <= xx_9;
    end
    if (reset) begin
      _T_584_4 <= 2'h0;
    end else begin
      _T_584_4 <= xx_15;
    end
    if (reset) begin
      _T_584_5 <= 2'h0;
    end else begin
      _T_584_5 <= xx_16;
    end
    if (reset) begin
      _T_584_7 <= 2'h0;
    end else begin
      _T_584_7 <= xx_22;
    end
    if (reset) begin
      _T_584_8 <= 2'h0;
    end else begin
      _T_584_8 <= xx_23;
    end
    if (reset) begin
      _T_661_1 <= 2'h0;
    end else begin
      _T_661_1 <= xx_15;
    end
    if (reset) begin
      _T_661_2 <= 2'h0;
    end else begin
      _T_661_2 <= xx_16;
    end
    if (reset) begin
      _T_661_4 <= 2'h0;
    end else begin
      _T_661_4 <= xx_22;
    end
    if (reset) begin
      _T_661_5 <= 2'h0;
    end else begin
      _T_661_5 <= xx_23;
    end
    if (reset) begin
      _T_661_7 <= 2'h0;
    end else begin
      _T_661_7 <= xx_29;
    end
    if (reset) begin
      _T_661_8 <= 2'h0;
    end else begin
      _T_661_8 <= xx_30;
    end
    if (reset) begin
      _T_738_1 <= 2'h0;
    end else begin
      _T_738_1 <= xx_22;
    end
    if (reset) begin
      _T_738_2 <= 2'h0;
    end else begin
      _T_738_2 <= xx_23;
    end
    if (reset) begin
      _T_738_4 <= 2'h0;
    end else begin
      _T_738_4 <= xx_29;
    end
    if (reset) begin
      _T_738_5 <= 2'h0;
    end else begin
      _T_738_5 <= xx_30;
    end
    if (reset) begin
      _T_738_7 <= 2'h0;
    end else begin
      _T_738_7 <= xx_36;
    end
    if (reset) begin
      _T_738_8 <= 2'h0;
    end else begin
      _T_738_8 <= xx_37;
    end
    if (reset) begin
      _T_815_1 <= 2'h0;
    end else begin
      _T_815_1 <= xx_29;
    end
    if (reset) begin
      _T_815_2 <= 2'h0;
    end else begin
      _T_815_2 <= xx_30;
    end
    if (reset) begin
      _T_815_4 <= 2'h0;
    end else begin
      _T_815_4 <= xx_36;
    end
    if (reset) begin
      _T_815_5 <= 2'h0;
    end else begin
      _T_815_5 <= xx_37;
    end
    if (reset) begin
      _T_892_3 <= 2'h0;
    end else begin
      _T_892_3 <= xx_8;
    end
    if (reset) begin
      _T_892_4 <= 2'h0;
    end else begin
      _T_892_4 <= xx_9;
    end
    if (reset) begin
      _T_892_5 <= 2'h0;
    end else begin
      _T_892_5 <= xx_10;
    end
    if (reset) begin
      _T_892_6 <= 2'h0;
    end else begin
      _T_892_6 <= xx_15;
    end
    if (reset) begin
      _T_892_7 <= 2'h0;
    end else begin
      _T_892_7 <= xx_16;
    end
    if (reset) begin
      _T_892_8 <= 2'h0;
    end else begin
      _T_892_8 <= xx_17;
    end
    if (reset) begin
      _T_969_0 <= 2'h0;
    end else begin
      _T_969_0 <= xx_8;
    end
    if (reset) begin
      _T_969_1 <= 2'h0;
    end else begin
      _T_969_1 <= xx_9;
    end
    if (reset) begin
      _T_969_2 <= 2'h0;
    end else begin
      _T_969_2 <= xx_10;
    end
    if (reset) begin
      _T_969_3 <= 2'h0;
    end else begin
      _T_969_3 <= xx_15;
    end
    if (reset) begin
      _T_969_4 <= 2'h0;
    end else begin
      _T_969_4 <= xx_16;
    end
    if (reset) begin
      _T_969_5 <= 2'h0;
    end else begin
      _T_969_5 <= xx_17;
    end
    if (reset) begin
      _T_969_6 <= 2'h0;
    end else begin
      _T_969_6 <= xx_22;
    end
    if (reset) begin
      _T_969_7 <= 2'h0;
    end else begin
      _T_969_7 <= xx_23;
    end
    if (reset) begin
      _T_969_8 <= 2'h0;
    end else begin
      _T_969_8 <= xx_24;
    end
    if (reset) begin
      _T_1046_0 <= 2'h0;
    end else begin
      _T_1046_0 <= xx_15;
    end
    if (reset) begin
      _T_1046_1 <= 2'h0;
    end else begin
      _T_1046_1 <= xx_16;
    end
    if (reset) begin
      _T_1046_2 <= 2'h0;
    end else begin
      _T_1046_2 <= xx_17;
    end
    if (reset) begin
      _T_1046_3 <= 2'h0;
    end else begin
      _T_1046_3 <= xx_22;
    end
    if (reset) begin
      _T_1046_4 <= 2'h0;
    end else begin
      _T_1046_4 <= xx_23;
    end
    if (reset) begin
      _T_1046_5 <= 2'h0;
    end else begin
      _T_1046_5 <= xx_24;
    end
    if (reset) begin
      _T_1046_6 <= 2'h0;
    end else begin
      _T_1046_6 <= xx_29;
    end
    if (reset) begin
      _T_1046_7 <= 2'h0;
    end else begin
      _T_1046_7 <= xx_30;
    end
    if (reset) begin
      _T_1046_8 <= 2'h0;
    end else begin
      _T_1046_8 <= xx_31;
    end
    if (reset) begin
      _T_1123_0 <= 2'h0;
    end else begin
      _T_1123_0 <= xx_22;
    end
    if (reset) begin
      _T_1123_1 <= 2'h0;
    end else begin
      _T_1123_1 <= xx_23;
    end
    if (reset) begin
      _T_1123_2 <= 2'h0;
    end else begin
      _T_1123_2 <= xx_24;
    end
    if (reset) begin
      _T_1123_3 <= 2'h0;
    end else begin
      _T_1123_3 <= xx_29;
    end
    if (reset) begin
      _T_1123_4 <= 2'h0;
    end else begin
      _T_1123_4 <= xx_30;
    end
    if (reset) begin
      _T_1123_5 <= 2'h0;
    end else begin
      _T_1123_5 <= xx_31;
    end
    if (reset) begin
      _T_1123_6 <= 2'h0;
    end else begin
      _T_1123_6 <= xx_36;
    end
    if (reset) begin
      _T_1123_7 <= 2'h0;
    end else begin
      _T_1123_7 <= xx_37;
    end
    if (reset) begin
      _T_1123_8 <= 2'h0;
    end else begin
      _T_1123_8 <= xx_38;
    end
    if (reset) begin
      _T_1200_0 <= 2'h0;
    end else begin
      _T_1200_0 <= xx_29;
    end
    if (reset) begin
      _T_1200_1 <= 2'h0;
    end else begin
      _T_1200_1 <= xx_30;
    end
    if (reset) begin
      _T_1200_2 <= 2'h0;
    end else begin
      _T_1200_2 <= xx_31;
    end
    if (reset) begin
      _T_1200_3 <= 2'h0;
    end else begin
      _T_1200_3 <= xx_36;
    end
    if (reset) begin
      _T_1200_4 <= 2'h0;
    end else begin
      _T_1200_4 <= xx_37;
    end
    if (reset) begin
      _T_1200_5 <= 2'h0;
    end else begin
      _T_1200_5 <= xx_38;
    end
    if (reset) begin
      _T_1277_3 <= 2'h0;
    end else begin
      _T_1277_3 <= xx_9;
    end
    if (reset) begin
      _T_1277_4 <= 2'h0;
    end else begin
      _T_1277_4 <= xx_10;
    end
    if (reset) begin
      _T_1277_5 <= 2'h0;
    end else begin
      _T_1277_5 <= xx_11;
    end
    if (reset) begin
      _T_1277_6 <= 2'h0;
    end else begin
      _T_1277_6 <= xx_16;
    end
    if (reset) begin
      _T_1277_7 <= 2'h0;
    end else begin
      _T_1277_7 <= xx_17;
    end
    if (reset) begin
      _T_1277_8 <= 2'h0;
    end else begin
      _T_1277_8 <= xx_18;
    end
    if (reset) begin
      _T_1354_0 <= 2'h0;
    end else begin
      _T_1354_0 <= xx_9;
    end
    if (reset) begin
      _T_1354_1 <= 2'h0;
    end else begin
      _T_1354_1 <= xx_10;
    end
    if (reset) begin
      _T_1354_2 <= 2'h0;
    end else begin
      _T_1354_2 <= xx_11;
    end
    if (reset) begin
      _T_1354_3 <= 2'h0;
    end else begin
      _T_1354_3 <= xx_16;
    end
    if (reset) begin
      _T_1354_4 <= 2'h0;
    end else begin
      _T_1354_4 <= xx_17;
    end
    if (reset) begin
      _T_1354_5 <= 2'h0;
    end else begin
      _T_1354_5 <= xx_18;
    end
    if (reset) begin
      _T_1354_6 <= 2'h0;
    end else begin
      _T_1354_6 <= xx_23;
    end
    if (reset) begin
      _T_1354_7 <= 2'h0;
    end else begin
      _T_1354_7 <= xx_24;
    end
    if (reset) begin
      _T_1354_8 <= 2'h0;
    end else begin
      _T_1354_8 <= xx_25;
    end
    if (reset) begin
      _T_1431_0 <= 2'h0;
    end else begin
      _T_1431_0 <= xx_16;
    end
    if (reset) begin
      _T_1431_1 <= 2'h0;
    end else begin
      _T_1431_1 <= xx_17;
    end
    if (reset) begin
      _T_1431_2 <= 2'h0;
    end else begin
      _T_1431_2 <= xx_18;
    end
    if (reset) begin
      _T_1431_3 <= 2'h0;
    end else begin
      _T_1431_3 <= xx_23;
    end
    if (reset) begin
      _T_1431_4 <= 2'h0;
    end else begin
      _T_1431_4 <= xx_24;
    end
    if (reset) begin
      _T_1431_5 <= 2'h0;
    end else begin
      _T_1431_5 <= xx_25;
    end
    if (reset) begin
      _T_1431_6 <= 2'h0;
    end else begin
      _T_1431_6 <= xx_30;
    end
    if (reset) begin
      _T_1431_7 <= 2'h0;
    end else begin
      _T_1431_7 <= xx_31;
    end
    if (reset) begin
      _T_1431_8 <= 2'h0;
    end else begin
      _T_1431_8 <= xx_32;
    end
    if (reset) begin
      _T_1508_0 <= 2'h0;
    end else begin
      _T_1508_0 <= xx_23;
    end
    if (reset) begin
      _T_1508_1 <= 2'h0;
    end else begin
      _T_1508_1 <= xx_24;
    end
    if (reset) begin
      _T_1508_2 <= 2'h0;
    end else begin
      _T_1508_2 <= xx_25;
    end
    if (reset) begin
      _T_1508_3 <= 2'h0;
    end else begin
      _T_1508_3 <= xx_30;
    end
    if (reset) begin
      _T_1508_4 <= 2'h0;
    end else begin
      _T_1508_4 <= xx_31;
    end
    if (reset) begin
      _T_1508_5 <= 2'h0;
    end else begin
      _T_1508_5 <= xx_32;
    end
    if (reset) begin
      _T_1508_6 <= 2'h0;
    end else begin
      _T_1508_6 <= xx_37;
    end
    if (reset) begin
      _T_1508_7 <= 2'h0;
    end else begin
      _T_1508_7 <= xx_38;
    end
    if (reset) begin
      _T_1508_8 <= 2'h0;
    end else begin
      _T_1508_8 <= xx_39;
    end
    if (reset) begin
      _T_1585_0 <= 2'h0;
    end else begin
      _T_1585_0 <= xx_30;
    end
    if (reset) begin
      _T_1585_1 <= 2'h0;
    end else begin
      _T_1585_1 <= xx_31;
    end
    if (reset) begin
      _T_1585_2 <= 2'h0;
    end else begin
      _T_1585_2 <= xx_32;
    end
    if (reset) begin
      _T_1585_3 <= 2'h0;
    end else begin
      _T_1585_3 <= xx_37;
    end
    if (reset) begin
      _T_1585_4 <= 2'h0;
    end else begin
      _T_1585_4 <= xx_38;
    end
    if (reset) begin
      _T_1585_5 <= 2'h0;
    end else begin
      _T_1585_5 <= xx_39;
    end
    if (reset) begin
      _T_1662_3 <= 2'h0;
    end else begin
      _T_1662_3 <= xx_10;
    end
    if (reset) begin
      _T_1662_4 <= 2'h0;
    end else begin
      _T_1662_4 <= xx_11;
    end
    if (reset) begin
      _T_1662_5 <= 2'h0;
    end else begin
      _T_1662_5 <= xx_12;
    end
    if (reset) begin
      _T_1662_6 <= 2'h0;
    end else begin
      _T_1662_6 <= xx_17;
    end
    if (reset) begin
      _T_1662_7 <= 2'h0;
    end else begin
      _T_1662_7 <= xx_18;
    end
    if (reset) begin
      _T_1662_8 <= 2'h0;
    end else begin
      _T_1662_8 <= xx_19;
    end
    if (reset) begin
      _T_1739_0 <= 2'h0;
    end else begin
      _T_1739_0 <= xx_10;
    end
    if (reset) begin
      _T_1739_1 <= 2'h0;
    end else begin
      _T_1739_1 <= xx_11;
    end
    if (reset) begin
      _T_1739_2 <= 2'h0;
    end else begin
      _T_1739_2 <= xx_12;
    end
    if (reset) begin
      _T_1739_3 <= 2'h0;
    end else begin
      _T_1739_3 <= xx_17;
    end
    if (reset) begin
      _T_1739_4 <= 2'h0;
    end else begin
      _T_1739_4 <= xx_18;
    end
    if (reset) begin
      _T_1739_5 <= 2'h0;
    end else begin
      _T_1739_5 <= xx_19;
    end
    if (reset) begin
      _T_1739_6 <= 2'h0;
    end else begin
      _T_1739_6 <= xx_24;
    end
    if (reset) begin
      _T_1739_7 <= 2'h0;
    end else begin
      _T_1739_7 <= xx_25;
    end
    if (reset) begin
      _T_1739_8 <= 2'h0;
    end else begin
      _T_1739_8 <= xx_26;
    end
    if (reset) begin
      _T_1816_0 <= 2'h0;
    end else begin
      _T_1816_0 <= xx_17;
    end
    if (reset) begin
      _T_1816_1 <= 2'h0;
    end else begin
      _T_1816_1 <= xx_18;
    end
    if (reset) begin
      _T_1816_2 <= 2'h0;
    end else begin
      _T_1816_2 <= xx_19;
    end
    if (reset) begin
      _T_1816_3 <= 2'h0;
    end else begin
      _T_1816_3 <= xx_24;
    end
    if (reset) begin
      _T_1816_4 <= 2'h0;
    end else begin
      _T_1816_4 <= xx_25;
    end
    if (reset) begin
      _T_1816_5 <= 2'h0;
    end else begin
      _T_1816_5 <= xx_26;
    end
    if (reset) begin
      _T_1816_6 <= 2'h0;
    end else begin
      _T_1816_6 <= xx_31;
    end
    if (reset) begin
      _T_1816_7 <= 2'h0;
    end else begin
      _T_1816_7 <= xx_32;
    end
    if (reset) begin
      _T_1816_8 <= 2'h0;
    end else begin
      _T_1816_8 <= xx_33;
    end
    if (reset) begin
      _T_1893_0 <= 2'h0;
    end else begin
      _T_1893_0 <= xx_24;
    end
    if (reset) begin
      _T_1893_1 <= 2'h0;
    end else begin
      _T_1893_1 <= xx_25;
    end
    if (reset) begin
      _T_1893_2 <= 2'h0;
    end else begin
      _T_1893_2 <= xx_26;
    end
    if (reset) begin
      _T_1893_3 <= 2'h0;
    end else begin
      _T_1893_3 <= xx_31;
    end
    if (reset) begin
      _T_1893_4 <= 2'h0;
    end else begin
      _T_1893_4 <= xx_32;
    end
    if (reset) begin
      _T_1893_5 <= 2'h0;
    end else begin
      _T_1893_5 <= xx_33;
    end
    if (reset) begin
      _T_1893_6 <= 2'h0;
    end else begin
      _T_1893_6 <= xx_38;
    end
    if (reset) begin
      _T_1893_7 <= 2'h0;
    end else begin
      _T_1893_7 <= xx_39;
    end
    if (reset) begin
      _T_1893_8 <= 2'h0;
    end else begin
      _T_1893_8 <= xx_40;
    end
    if (reset) begin
      _T_1970_0 <= 2'h0;
    end else begin
      _T_1970_0 <= xx_31;
    end
    if (reset) begin
      _T_1970_1 <= 2'h0;
    end else begin
      _T_1970_1 <= xx_32;
    end
    if (reset) begin
      _T_1970_2 <= 2'h0;
    end else begin
      _T_1970_2 <= xx_33;
    end
    if (reset) begin
      _T_1970_3 <= 2'h0;
    end else begin
      _T_1970_3 <= xx_38;
    end
    if (reset) begin
      _T_1970_4 <= 2'h0;
    end else begin
      _T_1970_4 <= xx_39;
    end
    if (reset) begin
      _T_1970_5 <= 2'h0;
    end else begin
      _T_1970_5 <= xx_40;
    end
    if (reset) begin
      _T_2047_3 <= 2'h0;
    end else begin
      _T_2047_3 <= xx_11;
    end
    if (reset) begin
      _T_2047_4 <= 2'h0;
    end else begin
      _T_2047_4 <= xx_12;
    end
    if (reset) begin
      _T_2047_6 <= 2'h0;
    end else begin
      _T_2047_6 <= xx_18;
    end
    if (reset) begin
      _T_2047_7 <= 2'h0;
    end else begin
      _T_2047_7 <= xx_19;
    end
    if (reset) begin
      _T_2124_0 <= 2'h0;
    end else begin
      _T_2124_0 <= xx_11;
    end
    if (reset) begin
      _T_2124_1 <= 2'h0;
    end else begin
      _T_2124_1 <= xx_12;
    end
    if (reset) begin
      _T_2124_3 <= 2'h0;
    end else begin
      _T_2124_3 <= xx_18;
    end
    if (reset) begin
      _T_2124_4 <= 2'h0;
    end else begin
      _T_2124_4 <= xx_19;
    end
    if (reset) begin
      _T_2124_6 <= 2'h0;
    end else begin
      _T_2124_6 <= xx_25;
    end
    if (reset) begin
      _T_2124_7 <= 2'h0;
    end else begin
      _T_2124_7 <= xx_26;
    end
    if (reset) begin
      _T_2201_0 <= 2'h0;
    end else begin
      _T_2201_0 <= xx_18;
    end
    if (reset) begin
      _T_2201_1 <= 2'h0;
    end else begin
      _T_2201_1 <= xx_19;
    end
    if (reset) begin
      _T_2201_3 <= 2'h0;
    end else begin
      _T_2201_3 <= xx_25;
    end
    if (reset) begin
      _T_2201_4 <= 2'h0;
    end else begin
      _T_2201_4 <= xx_26;
    end
    if (reset) begin
      _T_2201_6 <= 2'h0;
    end else begin
      _T_2201_6 <= xx_32;
    end
    if (reset) begin
      _T_2201_7 <= 2'h0;
    end else begin
      _T_2201_7 <= xx_33;
    end
    if (reset) begin
      _T_2278_0 <= 2'h0;
    end else begin
      _T_2278_0 <= xx_25;
    end
    if (reset) begin
      _T_2278_1 <= 2'h0;
    end else begin
      _T_2278_1 <= xx_26;
    end
    if (reset) begin
      _T_2278_3 <= 2'h0;
    end else begin
      _T_2278_3 <= xx_32;
    end
    if (reset) begin
      _T_2278_4 <= 2'h0;
    end else begin
      _T_2278_4 <= xx_33;
    end
    if (reset) begin
      _T_2278_6 <= 2'h0;
    end else begin
      _T_2278_6 <= xx_39;
    end
    if (reset) begin
      _T_2278_7 <= 2'h0;
    end else begin
      _T_2278_7 <= xx_40;
    end
    if (reset) begin
      _T_2355_0 <= 2'h0;
    end else begin
      _T_2355_0 <= xx_32;
    end
    if (reset) begin
      _T_2355_1 <= 2'h0;
    end else begin
      _T_2355_1 <= xx_33;
    end
    if (reset) begin
      _T_2355_3 <= 2'h0;
    end else begin
      _T_2355_3 <= xx_39;
    end
    if (reset) begin
      _T_2355_4 <= 2'h0;
    end else begin
      _T_2355_4 <= xx_40;
    end
  end
endmodule
